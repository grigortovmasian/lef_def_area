#----------------------------------------------------------------------------
# Description	: Cell LEF definitions for ts18ugfsdmp
#		  (TSMC 018um fsg -StdVt Metal Programable Library)
# Date		: $Date: 2006/06/08 03:58:23 $
# Copyright	: 1997-2006 by Virage Logic Corporation
# Revision	: Version $Revision: 1.18 $
#----------------------------------------------------------------------------

VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

# Placement site definition for this library.
SITE ts18_dmp
  CLASS core ;
  SIZE 2.24 BY 5.6 ;
END ts18_dmp

#----------------------------------------------------------------------------
# Cell macro definitions.
#-----------------------------------------------------------------------
#      Cell        : MDN_ADDF_1
#      Description : Full adder
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ADDF_1
  CLASS CORE ;
  FOREIGN MDN_ADDF_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.975 2.43 4.34 2.61 ;
      RECT  3.805 2.61 4.34 2.685 ;
      RECT  3.805 2.685 9.075 2.915 ;
      RECT  7.165 2.35 7.395 2.685 ;
      RECT  3.805 2.915 4.035 3.49 ;
      RECT  8.845 2.915 9.075 3.49 ;
      RECT  1.54 2.125 1.82 3.49 ;
      RECT  1.54 3.49 4.035 3.72 ;
      RECT  8.845 3.49 11.875 3.72 ;
      RECT  11.645 2.35 11.875 3.49 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 2.325 12.77 2.665 ;
      RECT  12.205 2.665 12.435 3.95 ;
      RECT  9.94 3.95 12.435 4.18 ;
      RECT  9.94 4.18 10.27 4.41 ;
      RECT  4.975 4.41 10.27 4.64 ;
      RECT  4.975 4.64 5.205 5.0 ;
      RECT  5.99 4.64 6.22 5.0 ;
      RECT  0.42 2.125 0.7 3.95 ;
      RECT  0.42 3.95 3.475 4.18 ;
      RECT  3.17 4.18 3.475 4.375 ;
      RECT  3.245 4.375 3.475 5.0 ;
      RECT  3.245 5.0 5.21 5.23 ;
      RECT  5.99 5.0 6.33 5.23 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.62 1.565 14.115 1.795 ;
      RECT  13.885 1.795 14.115 3.245 ;
      RECT  13.62 3.245 14.115 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 3.245 ;
      RECT  15.005 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.92 4.365 14.67 4.39 ;
      RECT  12.92 4.39 14.675 4.595 ;
      RECT  14.445 4.595 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.695 ;
      RECT  12.32 -0.14 12.995 0.14 ;
      RECT  12.765 0.14 12.995 1.005 ;
      RECT  12.765 1.005 13.26 1.235 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.52 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.52 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  9.965 0.37 10.81 0.6 ;
      RECT  9.965 0.6 10.195 0.76 ;
      RECT  2.61 0.37 3.475 0.6 ;
      RECT  3.245 0.6 3.475 0.76 ;
      RECT  3.245 0.76 10.195 0.99 ;
      RECT  8.23 0.37 8.57 0.76 ;
      RECT  0.14 1.005 2.76 1.235 ;
      RECT  10.63 1.005 11.72 1.235 ;
      RECT  3.915 1.22 5.0 1.45 ;
      RECT  6.15 1.22 9.48 1.45 ;
      RECT  9.91 1.565 13.24 1.795 ;
      RECT  9.91 1.795 10.14 3.03 ;
      RECT  13.01 1.795 13.24 3.805 ;
      RECT  9.91 3.03 10.25 3.26 ;
      RECT  13.01 3.805 15.18 4.035 ;
      RECT  14.95 4.035 15.18 5.0 ;
      RECT  14.95 5.0 15.29 5.23 ;
      RECT  3.245 1.68 9.635 1.91 ;
      RECT  9.405 1.91 9.635 2.7 ;
      RECT  3.245 1.91 3.475 3.03 ;
      RECT  3.19 3.03 3.53 3.26 ;
      RECT  6.2 3.805 8.515 3.95 ;
      RECT  6.2 3.95 9.48 4.035 ;
      RECT  8.285 4.035 9.48 4.18 ;
      RECT  4.365 3.805 5.0 4.035 ;
      RECT  4.365 4.035 4.595 4.365 ;
      RECT  3.91 4.365 4.595 4.595 ;
      RECT  0.18 4.41 2.76 4.64 ;
      RECT  10.63 4.42 11.72 4.65 ;
      RECT  9.35 5.0 14.17 5.23 ;
  END
END MDN_ADDF_1
#-----------------------------------------------------------------------
#      Cell        : MDN_ADDF_2
#      Description : Full adder
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ADDF_2
  CLASS CORE ;
  FOREIGN MDN_ADDF_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 2.35 4.035 2.66 ;
      RECT  3.805 2.66 9.07 2.685 ;
      RECT  7.165 2.35 7.395 2.66 ;
      RECT  3.805 2.685 9.075 2.94 ;
      RECT  3.805 2.94 4.035 3.49 ;
      RECT  8.845 2.94 9.075 3.49 ;
      RECT  1.54 2.125 1.82 3.49 ;
      RECT  1.54 3.49 4.035 3.72 ;
      RECT  8.845 3.49 11.875 3.72 ;
      RECT  11.645 2.35 11.875 3.49 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 2.43 12.905 2.66 ;
      RECT  12.205 2.66 12.435 3.95 ;
      RECT  9.94 3.95 12.435 4.18 ;
      RECT  9.94 4.18 10.27 4.41 ;
      RECT  4.98 4.41 10.27 4.64 ;
      RECT  4.98 4.64 5.21 5.0 ;
      RECT  5.99 4.64 6.22 5.0 ;
      RECT  0.42 2.125 0.7 3.95 ;
      RECT  0.42 3.95 3.5 4.18 ;
      RECT  3.17 4.18 3.5 4.34 ;
      RECT  3.22 4.34 3.5 5.0 ;
      RECT  3.22 5.0 5.21 5.23 ;
      RECT  5.99 5.0 6.33 5.23 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.62 1.565 15.795 1.795 ;
      RECT  15.565 1.795 15.795 3.245 ;
      RECT  13.62 3.245 15.795 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.86 1.005 16.355 1.235 ;
      RECT  16.125 1.235 16.355 1.565 ;
      RECT  16.125 1.565 17.74 1.795 ;
      RECT  16.685 1.795 16.915 3.245 ;
      RECT  16.125 3.245 17.755 3.475 ;
      RECT  16.125 3.475 16.355 3.805 ;
      RECT  15.86 3.805 16.355 4.035 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.87 4.365 14.675 4.595 ;
      RECT  14.445 4.595 14.675 5.46 ;
      RECT  14.445 5.46 18.09 5.74 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  7.725 4.905 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.905 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.905 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.695 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.695 ;
      RECT  12.32 -0.14 12.995 0.14 ;
      RECT  12.765 0.14 12.995 1.005 ;
      RECT  12.765 1.005 13.26 1.235 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.52 ;
      RECT  7.725 0.14 7.955 0.52 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  9.965 0.37 10.81 0.6 ;
      RECT  9.965 0.6 10.195 0.755 ;
      RECT  2.61 0.37 3.475 0.6 ;
      RECT  3.245 0.6 3.475 0.755 ;
      RECT  3.245 0.755 10.195 0.985 ;
      RECT  8.23 0.37 8.57 0.755 ;
      RECT  0.14 1.005 2.76 1.235 ;
      RECT  10.675 1.005 11.725 1.235 ;
      RECT  3.915 1.215 5.0 1.445 ;
      RECT  6.2 1.215 9.48 1.445 ;
      RECT  3.24 1.675 9.635 1.905 ;
      RECT  9.405 1.905 9.635 2.69 ;
      RECT  3.24 1.905 3.47 3.03 ;
      RECT  3.19 3.03 3.53 3.26 ;
      RECT  13.83 2.38 15.235 2.61 ;
      RECT  6.2 3.805 8.515 3.95 ;
      RECT  6.2 3.95 9.48 4.035 ;
      RECT  8.285 4.035 9.48 4.18 ;
      RECT  4.365 3.805 5.0 4.035 ;
      RECT  4.365 4.035 4.595 4.365 ;
      RECT  3.91 4.365 4.595 4.595 ;
      RECT  16.2 4.365 17.41 4.595 ;
      RECT  16.2 4.595 16.43 5.0 ;
      RECT  17.18 4.595 17.41 5.0 ;
      RECT  9.965 1.565 13.375 1.795 ;
      RECT  9.965 1.795 10.195 3.03 ;
      RECT  13.145 1.795 13.375 3.805 ;
      RECT  9.91 3.03 10.25 3.26 ;
      RECT  13.145 3.805 15.235 4.035 ;
      RECT  15.005 4.035 15.235 5.0 ;
      RECT  15.005 5.0 16.43 5.23 ;
      RECT  17.18 5.0 17.53 5.23 ;
      RECT  0.14 4.41 2.76 4.64 ;
      RECT  10.63 4.41 11.72 4.64 ;
      RECT  9.33 5.0 14.19 5.23 ;
  END
END MDN_ADDF_2
#-----------------------------------------------------------------------
#      Cell        : MDN_ADDF_4
#      Description : Full adder
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ADDF_4
  CLASS CORE ;
  FOREIGN MDN_ADDF_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 2.35 4.035 3.22 ;
      RECT  3.805 3.22 9.075 3.49 ;
      RECT  7.165 2.35 7.395 3.22 ;
      RECT  1.54 2.125 1.82 3.245 ;
      RECT  1.54 3.245 2.915 3.475 ;
      RECT  2.685 3.475 2.915 3.49 ;
      RECT  2.685 3.49 11.875 3.5 ;
      RECT  11.645 2.335 11.875 3.49 ;
      RECT  2.685 3.5 4.035 3.71 ;
      RECT  8.845 3.5 11.875 3.72 ;
      RECT  2.685 3.71 4.03 3.72 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.94 3.95 12.46 4.18 ;
      RECT  12.13 4.18 12.46 4.34 ;
      RECT  9.94 4.18 10.27 4.41 ;
      RECT  12.18 4.34 12.46 5.0 ;
      RECT  4.98 4.41 10.27 4.64 ;
      RECT  4.98 4.64 5.21 5.0 ;
      RECT  6.1 4.64 6.33 5.0 ;
      RECT  0.42 2.125 0.7 3.805 ;
      RECT  0.42 3.805 2.355 3.95 ;
      RECT  0.42 3.95 3.5 4.035 ;
      RECT  2.125 4.035 3.5 4.18 ;
      RECT  3.17 4.18 3.5 4.34 ;
      RECT  3.22 4.34 3.5 5.0 ;
      RECT  3.22 5.0 5.21 5.23 ;
      RECT  5.99 5.0 6.33 5.23 ;
      RECT  12.18 5.0 13.05 5.23 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.62 1.565 17.74 1.795 ;
      RECT  15.565 1.795 15.795 3.245 ;
      RECT  13.58 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.06 1.565 22.22 1.795 ;
      RECT  20.045 1.795 20.275 3.245 ;
      RECT  18.06 3.245 22.22 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.905 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.87 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  12.92 4.365 14.675 4.595 ;
      RECT  14.445 4.595 14.675 5.46 ;
      RECT  14.445 5.46 16.915 5.74 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  7.725 4.905 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.695 ;
      RECT  18.925 -0.14 19.6 0.14 ;
      RECT  18.925 0.14 19.155 0.695 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.695 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.695 ;
      RECT  12.32 -0.14 12.995 0.14 ;
      RECT  12.765 0.14 12.995 0.89 ;
      RECT  12.765 0.89 13.26 1.12 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.52 ;
      RECT  7.725 0.14 7.955 0.52 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  2.63 0.37 3.475 0.6 ;
      RECT  3.245 0.6 3.475 0.755 ;
      RECT  3.245 0.755 8.57 0.985 ;
      RECT  8.23 0.37 8.57 0.755 ;
      RECT  9.35 0.37 12.435 0.6 ;
      RECT  9.35 0.6 9.58 1.215 ;
      RECT  12.205 0.6 12.435 1.35 ;
      RECT  3.245 1.215 9.585 1.445 ;
      RECT  12.205 1.35 13.385 1.58 ;
      RECT  3.245 1.445 3.475 3.03 ;
      RECT  13.155 1.58 13.385 2.405 ;
      RECT  13.155 2.405 15.29 2.635 ;
      RECT  3.19 3.03 3.53 3.26 ;
      RECT  19.42 0.37 20.895 0.6 ;
      RECT  0.14 1.005 2.76 1.235 ;
      RECT  10.68 1.005 11.72 1.235 ;
      RECT  9.91 1.565 11.315 1.795 ;
      RECT  11.085 1.795 11.315 1.81 ;
      RECT  11.085 1.81 12.925 2.04 ;
      RECT  11.085 2.04 11.315 3.03 ;
      RECT  12.695 2.04 12.925 3.805 ;
      RECT  9.91 3.03 11.315 3.26 ;
      RECT  12.695 3.805 15.235 4.035 ;
      RECT  15.005 4.035 15.235 4.365 ;
      RECT  15.005 4.365 19.625 4.595 ;
      RECT  18.27 4.595 18.5 5.0 ;
      RECT  19.395 4.595 19.625 5.0 ;
      RECT  18.27 5.0 18.65 5.23 ;
      RECT  19.395 5.0 19.77 5.23 ;
      RECT  3.915 1.675 5.0 1.905 ;
      RECT  6.15 1.74 9.48 1.97 ;
      RECT  8.23 2.395 10.81 2.625 ;
      RECT  16.07 2.405 17.53 2.635 ;
      RECT  20.55 2.405 22.01 2.635 ;
      RECT  6.2 3.805 6.54 3.81 ;
      RECT  6.15 3.81 8.475 3.95 ;
      RECT  6.9 3.805 7.24 3.81 ;
      RECT  6.15 3.95 9.48 4.04 ;
      RECT  8.245 4.04 9.48 4.18 ;
      RECT  4.365 3.805 5.0 4.035 ;
      RECT  4.365 4.035 4.595 4.365 ;
      RECT  3.91 4.365 4.595 4.595 ;
      RECT  0.14 4.41 2.76 4.64 ;
      RECT  10.68 4.41 11.72 4.64 ;
      RECT  14.95 5.0 16.41 5.23 ;
  END
END MDN_ADDF_4
#-----------------------------------------------------------------------
#      Cell        : MDN_ADDF_P1_1
#      Description : Full adder
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ADDF_P1_1
  CLASS CORE ;
  FOREIGN MDN_ADDF_P1_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 2.35 4.035 3.5 ;
      RECT  3.17 3.5 4.035 3.56 ;
      RECT  1.54 2.125 1.82 3.5 ;
      RECT  1.54 3.5 1.87 3.56 ;
      RECT  1.54 3.56 4.035 3.79 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.245 1.565 17.74 1.795 ;
      RECT  17.245 1.795 17.475 3.245 ;
      RECT  17.245 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.86 1.565 16.915 1.795 ;
      RECT  16.685 1.795 16.915 3.245 ;
      RECT  15.86 3.245 16.915 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  12.205 5.08 12.435 5.46 ;
      RECT  11.76 5.46 12.88 5.74 ;
      RECT  9.965 5.08 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 5.08 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.805 4.48 4.3 4.71 ;
      RECT  3.805 4.71 4.035 5.46 ;
      RECT  3.805 5.46 4.48 5.74 ;
      RECT  1.005 5.08 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  12.205 -0.14 13.44 0.14 ;
      RECT  12.205 0.14 12.435 0.52 ;
      RECT  9.405 -0.14 10.08 0.14 ;
      RECT  9.405 0.14 9.635 0.89 ;
      RECT  9.14 0.89 9.635 1.12 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  12.765 0.37 15.29 0.6 ;
      RECT  12.765 0.6 12.995 0.825 ;
      RECT  9.965 0.825 12.995 1.055 ;
      RECT  9.965 1.055 10.195 1.4 ;
      RECT  5.99 0.37 7.185 0.6 ;
      RECT  6.955 0.6 7.185 1.29 ;
      RECT  6.955 1.29 8.985 1.295 ;
      RECT  6.955 1.295 8.99 1.3 ;
      RECT  6.955 1.3 8.995 1.305 ;
      RECT  6.955 1.305 9.0 1.31 ;
      RECT  6.955 1.31 9.005 1.315 ;
      RECT  6.955 1.315 9.01 1.32 ;
      RECT  6.955 1.32 9.015 1.325 ;
      RECT  6.955 1.325 9.02 1.33 ;
      RECT  6.955 1.33 9.025 1.335 ;
      RECT  6.955 1.335 9.03 1.34 ;
      RECT  6.955 1.34 9.035 1.345 ;
      RECT  6.955 1.345 9.04 1.35 ;
      RECT  6.955 1.35 9.045 1.355 ;
      RECT  6.955 1.355 9.05 1.36 ;
      RECT  6.955 1.36 9.055 1.365 ;
      RECT  6.955 1.365 9.06 1.37 ;
      RECT  6.955 1.37 9.065 1.375 ;
      RECT  6.955 1.375 9.07 1.38 ;
      RECT  6.955 1.38 9.075 1.385 ;
      RECT  6.955 1.385 9.08 1.39 ;
      RECT  6.955 1.39 9.085 1.395 ;
      RECT  6.955 1.395 9.09 1.4 ;
      RECT  6.955 1.4 10.195 1.52 ;
      RECT  8.88 1.52 10.195 1.525 ;
      RECT  6.955 1.52 7.395 1.535 ;
      RECT  8.885 1.525 10.195 1.53 ;
      RECT  8.89 1.53 10.195 1.535 ;
      RECT  7.165 1.535 7.395 3.03 ;
      RECT  8.895 1.535 10.195 1.54 ;
      RECT  8.9 1.54 10.195 1.545 ;
      RECT  8.905 1.545 10.195 1.55 ;
      RECT  8.91 1.55 10.195 1.555 ;
      RECT  8.915 1.555 10.195 1.56 ;
      RECT  8.92 1.56 10.195 1.565 ;
      RECT  8.925 1.565 10.195 1.57 ;
      RECT  8.93 1.57 10.195 1.575 ;
      RECT  8.935 1.575 10.195 1.58 ;
      RECT  8.94 1.58 10.195 1.585 ;
      RECT  8.945 1.585 10.195 1.59 ;
      RECT  8.95 1.59 10.195 1.595 ;
      RECT  8.955 1.595 10.195 1.6 ;
      RECT  8.96 1.6 10.195 1.605 ;
      RECT  8.965 1.605 10.195 1.61 ;
      RECT  8.97 1.61 10.195 1.615 ;
      RECT  8.975 1.615 10.195 1.62 ;
      RECT  8.98 1.62 10.195 1.625 ;
      RECT  8.985 1.625 10.195 1.63 ;
      RECT  6.9 3.03 7.395 3.26 ;
      RECT  4.065 0.83 6.705 1.005 ;
      RECT  1.005 1.005 6.705 1.06 ;
      RECT  6.2 1.06 6.705 1.12 ;
      RECT  1.005 1.06 4.295 1.235 ;
      RECT  6.475 1.12 6.705 2.1 ;
      RECT  1.005 1.235 1.235 4.02 ;
      RECT  6.475 2.1 6.855 2.38 ;
      RECT  0.18 4.02 5.0 4.25 ;
      RECT  14.435 1.005 15.5 1.01 ;
      RECT  14.43 1.01 15.5 1.015 ;
      RECT  14.425 1.015 15.5 1.02 ;
      RECT  14.42 1.02 15.5 1.025 ;
      RECT  14.415 1.025 15.5 1.03 ;
      RECT  14.41 1.03 15.5 1.035 ;
      RECT  14.405 1.035 15.5 1.04 ;
      RECT  14.4 1.04 15.5 1.045 ;
      RECT  14.395 1.045 15.5 1.05 ;
      RECT  14.39 1.05 15.5 1.055 ;
      RECT  14.385 1.055 15.5 1.06 ;
      RECT  14.38 1.06 15.5 1.065 ;
      RECT  14.375 1.065 15.5 1.07 ;
      RECT  14.37 1.07 15.5 1.075 ;
      RECT  14.365 1.075 15.5 1.08 ;
      RECT  14.36 1.08 15.5 1.085 ;
      RECT  14.355 1.085 15.5 1.09 ;
      RECT  14.35 1.09 15.5 1.095 ;
      RECT  14.345 1.095 15.5 1.1 ;
      RECT  14.34 1.1 15.5 1.105 ;
      RECT  14.335 1.105 15.5 1.11 ;
      RECT  14.33 1.11 15.5 1.115 ;
      RECT  14.325 1.115 15.5 1.12 ;
      RECT  14.32 1.12 15.5 1.125 ;
      RECT  14.315 1.125 15.5 1.13 ;
      RECT  14.31 1.13 15.5 1.135 ;
      RECT  14.305 1.135 15.5 1.14 ;
      RECT  14.3 1.14 15.5 1.145 ;
      RECT  14.295 1.145 15.5 1.15 ;
      RECT  14.29 1.15 15.5 1.155 ;
      RECT  14.285 1.155 15.5 1.16 ;
      RECT  14.28 1.16 15.5 1.165 ;
      RECT  14.275 1.165 15.5 1.17 ;
      RECT  14.27 1.17 15.5 1.175 ;
      RECT  14.265 1.175 15.5 1.18 ;
      RECT  14.26 1.18 15.5 1.185 ;
      RECT  14.255 1.185 15.5 1.19 ;
      RECT  14.25 1.19 15.5 1.195 ;
      RECT  14.245 1.195 15.5 1.2 ;
      RECT  14.24 1.2 15.5 1.205 ;
      RECT  14.235 1.205 15.5 1.21 ;
      RECT  14.23 1.21 15.5 1.215 ;
      RECT  14.225 1.215 15.5 1.22 ;
      RECT  14.22 1.22 15.5 1.225 ;
      RECT  14.215 1.225 15.5 1.23 ;
      RECT  14.21 1.23 15.5 1.235 ;
      RECT  14.205 1.235 14.53 1.24 ;
      RECT  14.2 1.24 14.525 1.245 ;
      RECT  14.195 1.245 14.52 1.25 ;
      RECT  14.19 1.25 14.515 1.255 ;
      RECT  14.185 1.255 14.51 1.26 ;
      RECT  14.18 1.26 14.505 1.265 ;
      RECT  14.175 1.265 14.5 1.27 ;
      RECT  14.17 1.27 14.495 1.275 ;
      RECT  14.165 1.275 14.49 1.28 ;
      RECT  14.16 1.28 14.485 1.285 ;
      RECT  14.155 1.285 14.48 1.29 ;
      RECT  14.15 1.29 14.475 1.295 ;
      RECT  14.145 1.295 14.47 1.3 ;
      RECT  14.14 1.3 14.465 1.305 ;
      RECT  14.135 1.305 14.46 1.31 ;
      RECT  14.13 1.31 14.455 1.315 ;
      RECT  14.125 1.315 14.45 1.32 ;
      RECT  14.12 1.32 14.445 1.325 ;
      RECT  14.115 1.325 14.44 1.33 ;
      RECT  14.11 1.33 14.435 1.335 ;
      RECT  14.105 1.335 14.43 1.34 ;
      RECT  14.1 1.34 14.425 1.345 ;
      RECT  14.095 1.345 14.42 1.35 ;
      RECT  14.09 1.35 14.415 1.355 ;
      RECT  14.085 1.355 14.41 1.36 ;
      RECT  14.08 1.36 14.405 1.365 ;
      RECT  14.075 1.365 14.4 1.37 ;
      RECT  14.07 1.37 14.395 1.375 ;
      RECT  14.065 1.375 14.39 1.38 ;
      RECT  14.06 1.38 14.385 1.385 ;
      RECT  14.055 1.385 14.38 1.39 ;
      RECT  14.05 1.39 14.375 1.395 ;
      RECT  14.045 1.395 14.37 1.4 ;
      RECT  14.04 1.4 14.365 1.405 ;
      RECT  14.035 1.405 14.36 1.41 ;
      RECT  14.03 1.41 14.355 1.415 ;
      RECT  14.025 1.415 14.35 1.42 ;
      RECT  14.02 1.42 14.345 1.425 ;
      RECT  14.015 1.425 14.34 1.43 ;
      RECT  14.01 1.43 14.335 1.435 ;
      RECT  14.005 1.435 14.33 1.44 ;
      RECT  14.0 1.44 14.325 1.445 ;
      RECT  13.995 1.445 14.32 1.45 ;
      RECT  13.99 1.45 14.315 1.455 ;
      RECT  13.985 1.455 14.31 1.46 ;
      RECT  13.98 1.46 14.305 1.465 ;
      RECT  13.975 1.465 14.3 1.47 ;
      RECT  13.97 1.47 14.295 1.475 ;
      RECT  13.965 1.475 14.29 1.48 ;
      RECT  13.96 1.48 14.285 1.485 ;
      RECT  13.955 1.485 14.28 1.49 ;
      RECT  13.95 1.49 14.275 1.495 ;
      RECT  13.945 1.495 14.27 1.5 ;
      RECT  13.94 1.5 14.265 1.505 ;
      RECT  13.935 1.505 14.26 1.51 ;
      RECT  13.93 1.51 14.255 1.515 ;
      RECT  13.925 1.515 14.25 1.52 ;
      RECT  13.92 1.52 14.245 1.525 ;
      RECT  13.915 1.525 14.24 1.53 ;
      RECT  13.91 1.53 14.235 1.535 ;
      RECT  13.905 1.535 14.23 1.54 ;
      RECT  13.9 1.54 14.225 1.545 ;
      RECT  13.895 1.545 14.22 1.55 ;
      RECT  13.89 1.55 14.215 1.555 ;
      RECT  13.885 1.555 14.21 1.56 ;
      RECT  13.88 1.56 14.205 1.565 ;
      RECT  13.875 1.565 14.2 1.57 ;
      RECT  13.87 1.57 14.195 1.575 ;
      RECT  13.865 1.575 14.19 1.58 ;
      RECT  13.86 1.58 14.185 1.585 ;
      RECT  13.855 1.585 14.18 1.59 ;
      RECT  13.85 1.59 14.175 1.595 ;
      RECT  13.845 1.595 14.17 1.6 ;
      RECT  13.84 1.6 14.165 1.605 ;
      RECT  13.835 1.605 14.16 1.61 ;
      RECT  13.83 1.61 14.155 1.615 ;
      RECT  13.825 1.615 14.15 1.62 ;
      RECT  13.82 1.62 14.145 1.625 ;
      RECT  13.815 1.625 14.14 1.63 ;
      RECT  13.81 1.63 14.135 1.635 ;
      RECT  13.805 1.635 14.13 1.64 ;
      RECT  13.8 1.64 14.125 1.645 ;
      RECT  13.795 1.645 14.12 1.65 ;
      RECT  13.79 1.65 14.115 1.655 ;
      RECT  13.785 1.655 14.11 1.66 ;
      RECT  13.78 1.66 14.105 1.665 ;
      RECT  13.775 1.665 14.1 1.67 ;
      RECT  13.77 1.67 14.095 1.675 ;
      RECT  13.765 1.675 14.09 1.68 ;
      RECT  13.76 1.68 14.085 1.685 ;
      RECT  13.755 1.685 14.08 1.69 ;
      RECT  13.75 1.69 14.075 1.695 ;
      RECT  13.745 1.695 14.07 1.7 ;
      RECT  13.74 1.7 14.065 1.705 ;
      RECT  13.735 1.705 14.06 1.71 ;
      RECT  13.73 1.71 14.055 1.715 ;
      RECT  13.725 1.715 14.05 1.72 ;
      RECT  13.72 1.72 14.045 1.725 ;
      RECT  13.715 1.725 14.04 1.73 ;
      RECT  13.71 1.73 14.035 1.735 ;
      RECT  13.705 1.735 14.03 1.74 ;
      RECT  13.7 1.74 14.025 1.745 ;
      RECT  13.695 1.745 14.02 1.75 ;
      RECT  12.92 1.75 14.015 1.755 ;
      RECT  12.92 1.755 14.01 1.76 ;
      RECT  12.92 1.76 14.005 1.765 ;
      RECT  12.92 1.765 14.0 1.77 ;
      RECT  12.92 1.77 13.995 1.775 ;
      RECT  12.92 1.775 13.99 1.78 ;
      RECT  12.92 1.78 13.985 1.785 ;
      RECT  12.92 1.785 13.98 1.79 ;
      RECT  12.92 1.79 13.975 1.795 ;
      RECT  12.92 1.795 13.97 1.8 ;
      RECT  12.92 1.8 13.965 1.805 ;
      RECT  12.92 1.805 13.96 1.81 ;
      RECT  12.92 1.81 13.955 1.815 ;
      RECT  12.92 1.815 13.95 1.82 ;
      RECT  12.92 1.82 13.945 1.825 ;
      RECT  12.92 1.825 13.94 1.83 ;
      RECT  12.92 1.83 13.935 1.835 ;
      RECT  12.92 1.835 13.93 1.84 ;
      RECT  12.92 1.84 13.925 1.845 ;
      RECT  12.92 1.845 13.92 1.85 ;
      RECT  12.92 1.85 13.915 1.855 ;
      RECT  12.92 1.855 13.91 1.86 ;
      RECT  12.92 1.86 13.905 1.865 ;
      RECT  12.92 1.865 13.9 1.87 ;
      RECT  12.92 1.87 13.895 1.875 ;
      RECT  12.92 1.875 13.89 1.88 ;
      RECT  12.92 1.88 13.885 1.885 ;
      RECT  12.92 1.885 13.88 1.89 ;
      RECT  12.92 1.89 13.875 1.895 ;
      RECT  12.92 1.895 13.87 1.9 ;
      RECT  12.92 1.9 13.865 1.905 ;
      RECT  12.92 1.905 13.86 1.91 ;
      RECT  12.92 1.91 13.855 1.915 ;
      RECT  12.92 1.915 13.85 1.92 ;
      RECT  12.92 1.92 13.845 1.925 ;
      RECT  12.92 1.925 13.84 1.93 ;
      RECT  12.92 1.93 13.835 1.935 ;
      RECT  12.92 1.935 13.83 1.94 ;
      RECT  12.92 1.94 13.825 1.945 ;
      RECT  12.92 1.945 13.82 1.95 ;
      RECT  12.92 1.95 13.815 1.955 ;
      RECT  12.92 1.955 13.81 1.96 ;
      RECT  12.92 1.96 13.805 1.965 ;
      RECT  12.92 1.965 13.8 1.97 ;
      RECT  12.92 1.97 13.795 1.975 ;
      RECT  12.92 1.975 13.79 1.98 ;
      RECT  13.325 1.98 13.555 3.24 ;
      RECT  12.92 3.24 13.96 3.47 ;
      RECT  13.325 0.89 13.96 1.12 ;
      RECT  13.325 1.12 13.555 1.29 ;
      RECT  11.38 1.29 13.555 1.52 ;
      RECT  12.205 1.52 12.435 2.435 ;
      RECT  12.205 2.435 13.05 2.665 ;
      RECT  12.205 2.665 12.435 3.245 ;
      RECT  11.37 3.245 12.435 3.475 ;
      RECT  12.205 3.475 12.435 3.7 ;
      RECT  12.205 3.7 15.5 3.93 ;
      RECT  10.68 1.565 11.075 1.795 ;
      RECT  10.845 1.795 11.075 2.41 ;
      RECT  10.845 2.41 11.93 2.64 ;
      RECT  10.845 2.64 11.075 3.245 ;
      RECT  9.14 3.245 11.075 3.475 ;
      RECT  5.43 1.75 5.77 1.98 ;
      RECT  5.485 1.98 5.715 4.16 ;
      RECT  5.485 4.16 14.675 4.365 ;
      RECT  5.485 4.365 17.42 4.39 ;
      RECT  14.445 4.39 17.42 4.595 ;
      RECT  17.19 4.595 17.42 5.0 ;
      RECT  17.19 5.0 17.53 5.23 ;
      RECT  8.44 1.75 8.78 1.98 ;
      RECT  8.55 1.98 8.78 2.445 ;
      RECT  8.55 2.445 9.69 2.675 ;
      RECT  8.55 2.675 8.78 3.245 ;
      RECT  8.44 3.245 8.78 3.475 ;
      RECT  14.39 1.75 14.73 1.98 ;
      RECT  14.445 1.98 14.675 2.445 ;
      RECT  14.445 2.445 16.41 2.675 ;
      RECT  14.445 2.675 14.675 3.455 ;
      RECT  9.955 2.1 10.595 2.38 ;
      RECT  10.365 2.38 10.595 2.68 ;
      RECT  8.06 2.36 8.29 2.685 ;
      RECT  7.725 2.685 8.29 2.915 ;
      RECT  7.725 2.915 7.955 3.615 ;
      RECT  4.77 1.29 5.975 1.295 ;
      RECT  4.77 1.295 5.98 1.3 ;
      RECT  4.77 1.3 5.985 1.305 ;
      RECT  4.77 1.305 5.99 1.31 ;
      RECT  4.77 1.31 5.995 1.315 ;
      RECT  4.77 1.315 6.0 1.32 ;
      RECT  4.77 1.32 6.005 1.325 ;
      RECT  4.77 1.325 6.01 1.33 ;
      RECT  4.77 1.33 6.015 1.335 ;
      RECT  4.77 1.335 6.02 1.34 ;
      RECT  4.77 1.34 6.025 1.345 ;
      RECT  4.77 1.345 6.03 1.35 ;
      RECT  4.77 1.35 6.035 1.355 ;
      RECT  4.77 1.355 6.04 1.36 ;
      RECT  4.77 1.36 6.045 1.365 ;
      RECT  4.77 1.365 6.05 1.37 ;
      RECT  4.77 1.37 6.055 1.375 ;
      RECT  4.77 1.375 6.06 1.38 ;
      RECT  4.77 1.38 6.065 1.385 ;
      RECT  4.77 1.385 6.07 1.39 ;
      RECT  4.77 1.39 6.075 1.395 ;
      RECT  4.77 1.395 6.08 1.4 ;
      RECT  4.77 1.4 6.085 1.405 ;
      RECT  4.77 1.405 6.09 1.41 ;
      RECT  4.77 1.41 6.095 1.415 ;
      RECT  4.77 1.415 6.1 1.42 ;
      RECT  4.77 1.42 6.105 1.425 ;
      RECT  4.77 1.425 6.11 1.43 ;
      RECT  4.77 1.43 6.115 1.435 ;
      RECT  4.77 1.435 6.12 1.44 ;
      RECT  4.77 1.44 6.125 1.445 ;
      RECT  4.77 1.445 6.13 1.45 ;
      RECT  4.77 1.45 6.135 1.455 ;
      RECT  4.77 1.455 6.14 1.46 ;
      RECT  4.77 1.46 6.145 1.465 ;
      RECT  4.77 1.465 6.15 1.47 ;
      RECT  4.77 1.47 6.155 1.475 ;
      RECT  4.77 1.475 6.16 1.48 ;
      RECT  4.77 1.48 6.165 1.485 ;
      RECT  4.77 1.485 6.17 1.49 ;
      RECT  4.77 1.49 6.175 1.495 ;
      RECT  4.77 1.495 6.18 1.5 ;
      RECT  4.77 1.5 6.185 1.505 ;
      RECT  4.77 1.505 6.19 1.51 ;
      RECT  4.77 1.51 6.195 1.515 ;
      RECT  4.77 1.515 6.2 1.52 ;
      RECT  5.87 1.52 6.205 1.525 ;
      RECT  4.77 1.52 5.0 1.565 ;
      RECT  5.875 1.525 6.21 1.53 ;
      RECT  5.88 1.53 6.215 1.535 ;
      RECT  5.885 1.535 6.22 1.54 ;
      RECT  5.89 1.54 6.225 1.545 ;
      RECT  5.895 1.545 6.23 1.55 ;
      RECT  5.9 1.55 6.23 1.555 ;
      RECT  5.905 1.555 6.23 1.56 ;
      RECT  5.91 1.56 6.23 1.565 ;
      RECT  2.42 1.565 5.0 1.795 ;
      RECT  5.915 1.565 6.23 1.57 ;
      RECT  5.92 1.57 6.23 1.575 ;
      RECT  5.925 1.575 6.23 1.58 ;
      RECT  5.93 1.58 6.23 1.585 ;
      RECT  5.935 1.585 6.23 1.59 ;
      RECT  5.94 1.59 6.23 1.595 ;
      RECT  5.945 1.595 6.23 1.6 ;
      RECT  5.95 1.6 6.23 1.605 ;
      RECT  5.955 1.605 6.23 1.61 ;
      RECT  5.96 1.61 6.23 1.615 ;
      RECT  5.965 1.615 6.23 1.62 ;
      RECT  5.97 1.62 6.23 1.625 ;
      RECT  5.975 1.625 6.23 1.63 ;
      RECT  5.98 1.63 6.23 1.635 ;
      RECT  5.985 1.635 6.23 1.64 ;
      RECT  5.99 1.64 6.23 1.645 ;
      RECT  5.995 1.645 6.23 1.65 ;
      RECT  6.0 1.65 6.23 3.615 ;
      RECT  2.685 1.795 2.915 3.1 ;
      RECT  2.42 3.1 2.915 3.33 ;
      RECT  6.0 3.615 7.955 3.845 ;
      RECT  0.5 4.62 1.72 4.85 ;
      RECT  1.49 4.85 1.72 4.925 ;
      RECT  0.5 4.85 0.73 5.0 ;
      RECT  1.49 4.925 2.97 5.155 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  2.43 5.155 2.97 5.18 ;
      RECT  2.63 5.18 2.97 5.23 ;
      RECT  7.22 4.62 14.06 4.85 ;
      RECT  13.81 4.85 14.06 4.9 ;
      RECT  7.22 4.85 7.45 5.0 ;
      RECT  13.83 4.9 14.06 5.0 ;
      RECT  4.87 5.0 7.45 5.23 ;
      RECT  13.83 5.0 14.17 5.23 ;
      LAYER METAL2 ;
      RECT  6.475 2.1 10.63 2.38 ;
      LAYER VIA12 ;
      RECT  6.535 2.11 6.795 2.37 ;
      RECT  10.015 2.11 10.275 2.37 ;
  END
END MDN_ADDF_P1_1
#-----------------------------------------------------------------------
#      Cell        : MDN_ADDF_P1_2
#      Description : Full adder
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ADDF_P1_2
  CLASS CORE ;
  FOREIGN MDN_ADDF_P1_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 3.495 ;
      RECT  1.54 3.495 4.035 3.725 ;
      RECT  3.805 2.35 4.035 3.495 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.1 1.565 19.98 1.795 ;
      RECT  18.925 1.795 19.155 3.245 ;
      RECT  18.1 3.245 19.98 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.86 1.565 17.74 1.795 ;
      RECT  16.685 1.795 16.915 3.245 ;
      RECT  15.86 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.87 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  12.15 5.135 12.49 5.46 ;
      RECT  11.76 5.46 12.88 5.74 ;
      RECT  9.965 4.875 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.875 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.805 4.415 4.3 4.645 ;
      RECT  3.805 4.645 4.035 5.46 ;
      RECT  3.805 5.46 4.65 5.74 ;
      RECT  1.005 4.95 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  15.51 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.595 ;
      RECT  9.405 -0.14 10.08 0.14 ;
      RECT  9.405 0.14 9.635 0.89 ;
      RECT  9.14 0.89 9.635 1.12 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  12.765 0.37 15.29 0.6 ;
      RECT  12.765 0.6 12.995 0.825 ;
      RECT  9.965 0.825 12.995 1.055 ;
      RECT  9.965 1.055 10.195 1.405 ;
      RECT  5.99 0.37 7.46 0.6 ;
      RECT  7.23 0.6 7.46 1.005 ;
      RECT  6.9 1.005 8.7 1.01 ;
      RECT  6.9 1.01 8.705 1.015 ;
      RECT  6.9 1.015 8.71 1.02 ;
      RECT  6.9 1.02 8.715 1.025 ;
      RECT  6.9 1.025 8.72 1.03 ;
      RECT  6.9 1.03 8.725 1.035 ;
      RECT  6.9 1.035 8.73 1.04 ;
      RECT  6.9 1.04 8.735 1.045 ;
      RECT  6.9 1.045 8.74 1.05 ;
      RECT  6.9 1.05 8.745 1.055 ;
      RECT  6.9 1.055 8.75 1.06 ;
      RECT  6.9 1.06 8.755 1.065 ;
      RECT  6.9 1.065 8.76 1.07 ;
      RECT  6.9 1.07 8.765 1.075 ;
      RECT  6.9 1.075 8.77 1.08 ;
      RECT  6.9 1.08 8.775 1.085 ;
      RECT  6.9 1.085 8.78 1.09 ;
      RECT  6.9 1.09 8.785 1.095 ;
      RECT  6.9 1.095 8.79 1.1 ;
      RECT  6.9 1.1 8.795 1.105 ;
      RECT  6.9 1.105 8.8 1.11 ;
      RECT  6.9 1.11 8.805 1.115 ;
      RECT  6.9 1.115 8.81 1.12 ;
      RECT  6.9 1.12 8.815 1.125 ;
      RECT  6.9 1.125 8.82 1.13 ;
      RECT  6.9 1.13 8.825 1.135 ;
      RECT  6.9 1.135 8.83 1.14 ;
      RECT  6.9 1.14 8.835 1.145 ;
      RECT  6.9 1.145 8.84 1.15 ;
      RECT  6.9 1.15 8.845 1.155 ;
      RECT  6.9 1.155 8.85 1.16 ;
      RECT  6.9 1.16 8.855 1.165 ;
      RECT  6.9 1.165 8.86 1.17 ;
      RECT  6.9 1.17 8.865 1.175 ;
      RECT  6.9 1.175 8.87 1.18 ;
      RECT  6.9 1.18 8.875 1.185 ;
      RECT  6.9 1.185 8.88 1.19 ;
      RECT  6.9 1.19 8.885 1.195 ;
      RECT  6.9 1.195 8.89 1.2 ;
      RECT  6.9 1.2 8.895 1.205 ;
      RECT  6.9 1.205 8.9 1.21 ;
      RECT  6.9 1.21 8.905 1.215 ;
      RECT  6.9 1.215 8.91 1.22 ;
      RECT  6.9 1.22 8.915 1.225 ;
      RECT  6.9 1.225 8.92 1.23 ;
      RECT  6.9 1.23 8.925 1.235 ;
      RECT  8.595 1.235 8.93 1.24 ;
      RECT  7.23 1.235 7.46 3.035 ;
      RECT  8.6 1.24 8.935 1.245 ;
      RECT  8.605 1.245 8.94 1.25 ;
      RECT  8.61 1.25 8.945 1.255 ;
      RECT  8.615 1.255 8.95 1.26 ;
      RECT  8.62 1.26 8.955 1.265 ;
      RECT  8.625 1.265 8.96 1.27 ;
      RECT  8.63 1.27 8.965 1.275 ;
      RECT  8.635 1.275 8.97 1.28 ;
      RECT  8.64 1.28 8.975 1.285 ;
      RECT  8.645 1.285 8.98 1.29 ;
      RECT  8.65 1.29 8.985 1.295 ;
      RECT  8.655 1.295 8.99 1.3 ;
      RECT  8.66 1.3 8.995 1.305 ;
      RECT  8.665 1.305 9.0 1.31 ;
      RECT  8.67 1.31 9.005 1.315 ;
      RECT  8.675 1.315 9.01 1.32 ;
      RECT  8.68 1.32 9.015 1.325 ;
      RECT  8.685 1.325 9.02 1.33 ;
      RECT  8.69 1.33 9.025 1.335 ;
      RECT  8.695 1.335 9.03 1.34 ;
      RECT  8.7 1.34 9.035 1.345 ;
      RECT  8.705 1.345 9.04 1.35 ;
      RECT  8.71 1.35 9.045 1.355 ;
      RECT  8.715 1.355 9.05 1.36 ;
      RECT  8.72 1.36 9.055 1.365 ;
      RECT  8.725 1.365 9.06 1.37 ;
      RECT  8.73 1.37 9.065 1.375 ;
      RECT  8.735 1.375 9.07 1.38 ;
      RECT  8.74 1.38 9.075 1.385 ;
      RECT  8.745 1.385 9.08 1.39 ;
      RECT  8.75 1.39 9.085 1.395 ;
      RECT  8.755 1.395 9.09 1.4 ;
      RECT  8.76 1.4 9.095 1.405 ;
      RECT  8.765 1.405 10.195 1.41 ;
      RECT  8.77 1.41 10.195 1.415 ;
      RECT  8.775 1.415 10.195 1.42 ;
      RECT  8.78 1.42 10.195 1.425 ;
      RECT  8.785 1.425 10.195 1.43 ;
      RECT  8.79 1.43 10.195 1.435 ;
      RECT  8.795 1.435 10.195 1.44 ;
      RECT  8.8 1.44 10.195 1.445 ;
      RECT  8.805 1.445 10.195 1.45 ;
      RECT  8.81 1.45 10.195 1.455 ;
      RECT  8.815 1.455 10.195 1.46 ;
      RECT  8.82 1.46 10.195 1.465 ;
      RECT  8.825 1.465 10.195 1.47 ;
      RECT  8.83 1.47 10.195 1.475 ;
      RECT  8.835 1.475 10.195 1.48 ;
      RECT  8.84 1.48 10.195 1.485 ;
      RECT  8.845 1.485 10.195 1.49 ;
      RECT  8.85 1.49 10.195 1.495 ;
      RECT  8.855 1.495 10.195 1.5 ;
      RECT  8.86 1.5 10.195 1.505 ;
      RECT  8.865 1.505 10.195 1.51 ;
      RECT  8.87 1.51 10.195 1.515 ;
      RECT  8.875 1.515 10.195 1.52 ;
      RECT  8.88 1.52 10.195 1.525 ;
      RECT  8.885 1.525 10.195 1.53 ;
      RECT  8.89 1.53 10.195 1.535 ;
      RECT  8.895 1.535 10.195 1.54 ;
      RECT  8.9 1.54 10.195 1.545 ;
      RECT  8.905 1.545 10.195 1.55 ;
      RECT  8.91 1.55 10.195 1.555 ;
      RECT  8.915 1.555 10.195 1.56 ;
      RECT  8.92 1.56 10.195 1.565 ;
      RECT  8.925 1.565 10.195 1.57 ;
      RECT  8.93 1.57 10.195 1.575 ;
      RECT  8.935 1.575 10.195 1.58 ;
      RECT  8.94 1.58 10.195 1.585 ;
      RECT  8.945 1.585 10.195 1.59 ;
      RECT  8.95 1.59 10.195 1.595 ;
      RECT  8.955 1.595 10.195 1.6 ;
      RECT  8.96 1.6 10.195 1.605 ;
      RECT  8.965 1.605 10.195 1.61 ;
      RECT  8.97 1.61 10.195 1.615 ;
      RECT  8.975 1.615 10.195 1.62 ;
      RECT  8.98 1.62 10.195 1.625 ;
      RECT  8.985 1.625 10.195 1.63 ;
      RECT  8.99 1.63 10.195 1.635 ;
      RECT  6.9 3.035 7.46 3.265 ;
      RECT  17.19 0.37 17.53 0.6 ;
      RECT  17.19 0.6 17.42 1.005 ;
      RECT  16.07 0.37 16.41 0.6 ;
      RECT  16.18 0.6 16.41 1.005 ;
      RECT  16.18 1.005 17.42 1.235 ;
      RECT  14.415 1.005 15.5 1.01 ;
      RECT  14.41 1.01 15.5 1.015 ;
      RECT  14.405 1.015 15.5 1.02 ;
      RECT  14.4 1.02 15.5 1.025 ;
      RECT  14.395 1.025 15.5 1.03 ;
      RECT  14.39 1.03 15.5 1.035 ;
      RECT  14.385 1.035 15.5 1.04 ;
      RECT  14.38 1.04 15.5 1.045 ;
      RECT  14.375 1.045 15.5 1.05 ;
      RECT  14.37 1.05 15.5 1.055 ;
      RECT  14.365 1.055 15.5 1.06 ;
      RECT  14.36 1.06 15.5 1.065 ;
      RECT  14.355 1.065 15.5 1.07 ;
      RECT  14.35 1.07 15.5 1.075 ;
      RECT  14.345 1.075 15.5 1.08 ;
      RECT  14.34 1.08 15.5 1.085 ;
      RECT  14.335 1.085 15.5 1.09 ;
      RECT  14.33 1.09 15.5 1.095 ;
      RECT  14.325 1.095 15.5 1.1 ;
      RECT  14.32 1.1 15.5 1.105 ;
      RECT  14.315 1.105 15.5 1.11 ;
      RECT  14.31 1.11 15.5 1.115 ;
      RECT  14.305 1.115 15.5 1.12 ;
      RECT  14.3 1.12 15.5 1.125 ;
      RECT  14.295 1.125 15.5 1.13 ;
      RECT  14.29 1.13 15.5 1.135 ;
      RECT  14.285 1.135 15.5 1.14 ;
      RECT  14.28 1.14 15.5 1.145 ;
      RECT  14.275 1.145 15.5 1.15 ;
      RECT  14.27 1.15 15.5 1.155 ;
      RECT  14.265 1.155 15.5 1.16 ;
      RECT  14.26 1.16 15.5 1.165 ;
      RECT  14.255 1.165 15.5 1.17 ;
      RECT  14.25 1.17 15.5 1.175 ;
      RECT  14.245 1.175 15.5 1.18 ;
      RECT  14.24 1.18 15.5 1.185 ;
      RECT  14.235 1.185 15.5 1.19 ;
      RECT  14.23 1.19 15.5 1.195 ;
      RECT  14.225 1.195 15.5 1.2 ;
      RECT  14.22 1.2 15.5 1.205 ;
      RECT  14.215 1.205 15.5 1.21 ;
      RECT  14.21 1.21 15.5 1.215 ;
      RECT  14.205 1.215 15.5 1.22 ;
      RECT  14.2 1.22 15.5 1.225 ;
      RECT  14.195 1.225 15.5 1.23 ;
      RECT  14.19 1.23 15.5 1.235 ;
      RECT  14.185 1.235 14.51 1.24 ;
      RECT  14.18 1.24 14.505 1.245 ;
      RECT  14.175 1.245 14.5 1.25 ;
      RECT  14.17 1.25 14.495 1.255 ;
      RECT  14.165 1.255 14.49 1.26 ;
      RECT  14.16 1.26 14.485 1.265 ;
      RECT  14.155 1.265 14.48 1.27 ;
      RECT  14.15 1.27 14.475 1.275 ;
      RECT  14.145 1.275 14.47 1.28 ;
      RECT  14.14 1.28 14.465 1.285 ;
      RECT  14.135 1.285 14.46 1.29 ;
      RECT  14.13 1.29 14.455 1.295 ;
      RECT  14.125 1.295 14.45 1.3 ;
      RECT  14.12 1.3 14.445 1.305 ;
      RECT  14.115 1.305 14.44 1.31 ;
      RECT  14.11 1.31 14.435 1.315 ;
      RECT  14.105 1.315 14.43 1.32 ;
      RECT  14.1 1.32 14.425 1.325 ;
      RECT  14.095 1.325 14.42 1.33 ;
      RECT  14.09 1.33 14.415 1.335 ;
      RECT  14.085 1.335 14.41 1.34 ;
      RECT  14.08 1.34 14.405 1.345 ;
      RECT  14.075 1.345 14.4 1.35 ;
      RECT  14.07 1.35 14.395 1.355 ;
      RECT  14.065 1.355 14.39 1.36 ;
      RECT  14.06 1.36 14.385 1.365 ;
      RECT  14.055 1.365 14.38 1.37 ;
      RECT  14.05 1.37 14.375 1.375 ;
      RECT  14.045 1.375 14.37 1.38 ;
      RECT  14.04 1.38 14.365 1.385 ;
      RECT  14.035 1.385 14.36 1.39 ;
      RECT  14.03 1.39 14.355 1.395 ;
      RECT  14.025 1.395 14.35 1.4 ;
      RECT  14.02 1.4 14.345 1.405 ;
      RECT  14.015 1.405 14.34 1.41 ;
      RECT  14.01 1.41 14.335 1.415 ;
      RECT  14.005 1.415 14.33 1.42 ;
      RECT  14.0 1.42 14.325 1.425 ;
      RECT  13.995 1.425 14.32 1.43 ;
      RECT  13.99 1.43 14.315 1.435 ;
      RECT  13.985 1.435 14.31 1.44 ;
      RECT  13.98 1.44 14.305 1.445 ;
      RECT  13.975 1.445 14.3 1.45 ;
      RECT  13.97 1.45 14.295 1.455 ;
      RECT  13.965 1.455 14.29 1.46 ;
      RECT  13.96 1.46 14.285 1.465 ;
      RECT  13.955 1.465 14.28 1.47 ;
      RECT  13.95 1.47 14.275 1.475 ;
      RECT  13.945 1.475 14.27 1.48 ;
      RECT  13.94 1.48 14.265 1.485 ;
      RECT  13.935 1.485 14.26 1.49 ;
      RECT  13.93 1.49 14.255 1.495 ;
      RECT  13.925 1.495 14.25 1.5 ;
      RECT  13.92 1.5 14.245 1.505 ;
      RECT  13.915 1.505 14.24 1.51 ;
      RECT  13.91 1.51 14.235 1.515 ;
      RECT  13.905 1.515 14.23 1.52 ;
      RECT  13.9 1.52 14.225 1.525 ;
      RECT  13.895 1.525 14.22 1.53 ;
      RECT  13.89 1.53 14.215 1.535 ;
      RECT  13.885 1.535 14.21 1.54 ;
      RECT  13.88 1.54 14.205 1.545 ;
      RECT  13.875 1.545 14.2 1.55 ;
      RECT  13.87 1.55 14.195 1.555 ;
      RECT  13.865 1.555 14.19 1.56 ;
      RECT  13.86 1.56 14.185 1.565 ;
      RECT  13.855 1.565 14.18 1.57 ;
      RECT  13.85 1.57 14.175 1.575 ;
      RECT  13.845 1.575 14.17 1.58 ;
      RECT  13.84 1.58 14.165 1.585 ;
      RECT  13.835 1.585 14.16 1.59 ;
      RECT  13.83 1.59 14.155 1.595 ;
      RECT  13.825 1.595 14.15 1.6 ;
      RECT  13.82 1.6 14.145 1.605 ;
      RECT  13.815 1.605 14.14 1.61 ;
      RECT  13.81 1.61 14.135 1.615 ;
      RECT  13.805 1.615 14.13 1.62 ;
      RECT  13.8 1.62 14.125 1.625 ;
      RECT  13.795 1.625 14.12 1.63 ;
      RECT  13.79 1.63 14.115 1.635 ;
      RECT  13.785 1.635 14.11 1.64 ;
      RECT  13.78 1.64 14.105 1.645 ;
      RECT  13.775 1.645 14.1 1.65 ;
      RECT  13.77 1.65 14.095 1.655 ;
      RECT  13.765 1.655 14.09 1.66 ;
      RECT  13.76 1.66 14.085 1.665 ;
      RECT  13.755 1.665 14.08 1.67 ;
      RECT  13.75 1.67 14.075 1.675 ;
      RECT  13.745 1.675 14.07 1.68 ;
      RECT  13.74 1.68 14.065 1.685 ;
      RECT  13.735 1.685 14.06 1.69 ;
      RECT  13.73 1.69 14.055 1.695 ;
      RECT  13.725 1.695 14.05 1.7 ;
      RECT  13.72 1.7 14.045 1.705 ;
      RECT  13.715 1.705 14.04 1.71 ;
      RECT  13.71 1.71 14.035 1.715 ;
      RECT  13.705 1.715 14.03 1.72 ;
      RECT  13.7 1.72 14.025 1.725 ;
      RECT  13.695 1.725 14.02 1.73 ;
      RECT  13.69 1.73 14.015 1.735 ;
      RECT  13.685 1.735 14.01 1.74 ;
      RECT  13.68 1.74 14.005 1.745 ;
      RECT  13.675 1.745 14.0 1.75 ;
      RECT  12.92 1.75 13.995 1.755 ;
      RECT  12.92 1.755 13.99 1.76 ;
      RECT  12.92 1.76 13.985 1.765 ;
      RECT  12.92 1.765 13.98 1.77 ;
      RECT  12.92 1.77 13.975 1.775 ;
      RECT  12.92 1.775 13.97 1.78 ;
      RECT  12.92 1.78 13.965 1.785 ;
      RECT  12.92 1.785 13.96 1.79 ;
      RECT  12.92 1.79 13.955 1.795 ;
      RECT  12.92 1.795 13.95 1.8 ;
      RECT  12.92 1.8 13.945 1.805 ;
      RECT  12.92 1.805 13.94 1.81 ;
      RECT  12.92 1.81 13.935 1.815 ;
      RECT  12.92 1.815 13.93 1.82 ;
      RECT  12.92 1.82 13.925 1.825 ;
      RECT  12.92 1.825 13.92 1.83 ;
      RECT  12.92 1.83 13.915 1.835 ;
      RECT  12.92 1.835 13.91 1.84 ;
      RECT  12.92 1.84 13.905 1.845 ;
      RECT  12.92 1.845 13.9 1.85 ;
      RECT  12.92 1.85 13.895 1.855 ;
      RECT  12.92 1.855 13.89 1.86 ;
      RECT  12.92 1.86 13.885 1.865 ;
      RECT  12.92 1.865 13.88 1.87 ;
      RECT  12.92 1.87 13.875 1.875 ;
      RECT  12.92 1.875 13.87 1.88 ;
      RECT  12.92 1.88 13.865 1.885 ;
      RECT  12.92 1.885 13.86 1.89 ;
      RECT  12.92 1.89 13.855 1.895 ;
      RECT  12.92 1.895 13.85 1.9 ;
      RECT  12.92 1.9 13.845 1.905 ;
      RECT  12.92 1.905 13.84 1.91 ;
      RECT  12.92 1.91 13.835 1.915 ;
      RECT  12.92 1.915 13.83 1.92 ;
      RECT  12.92 1.92 13.825 1.925 ;
      RECT  12.92 1.925 13.82 1.93 ;
      RECT  12.92 1.93 13.815 1.935 ;
      RECT  12.92 1.935 13.81 1.94 ;
      RECT  12.92 1.94 13.805 1.945 ;
      RECT  12.92 1.945 13.8 1.95 ;
      RECT  12.92 1.95 13.795 1.955 ;
      RECT  12.92 1.955 13.79 1.96 ;
      RECT  12.92 1.96 13.785 1.965 ;
      RECT  12.92 1.965 13.78 1.97 ;
      RECT  12.92 1.97 13.775 1.975 ;
      RECT  12.92 1.975 13.77 1.98 ;
      RECT  13.325 1.98 13.555 3.245 ;
      RECT  12.92 3.245 13.96 3.475 ;
      RECT  13.325 0.89 13.96 1.12 ;
      RECT  13.325 1.12 13.555 1.29 ;
      RECT  11.435 1.29 13.555 1.52 ;
      RECT  11.435 1.52 11.665 1.63 ;
      RECT  12.2 1.52 12.43 2.39 ;
      RECT  12.2 2.39 13.05 2.62 ;
      RECT  12.2 2.62 12.43 3.3 ;
      RECT  11.435 3.19 11.665 3.3 ;
      RECT  11.435 3.3 12.43 3.53 ;
      RECT  12.2 3.53 12.43 3.755 ;
      RECT  12.2 3.755 15.5 3.985 ;
      RECT  10.68 1.565 11.205 1.795 ;
      RECT  10.975 1.795 11.205 2.39 ;
      RECT  10.975 2.39 11.93 2.62 ;
      RECT  10.975 2.62 11.205 3.245 ;
      RECT  9.14 3.245 11.205 3.475 ;
      RECT  5.38 1.75 5.72 1.98 ;
      RECT  5.485 1.98 5.715 3.955 ;
      RECT  5.485 3.955 11.875 4.185 ;
      RECT  11.645 4.185 11.875 4.215 ;
      RECT  11.645 4.215 14.65 4.365 ;
      RECT  11.645 4.365 19.66 4.445 ;
      RECT  14.42 4.445 19.66 4.595 ;
      RECT  18.42 4.595 18.65 5.0 ;
      RECT  19.43 4.595 19.66 5.0 ;
      RECT  18.31 5.0 18.65 5.23 ;
      RECT  19.43 5.0 19.77 5.23 ;
      RECT  8.44 1.75 8.78 1.98 ;
      RECT  8.55 1.98 8.78 2.39 ;
      RECT  8.55 2.39 9.69 2.62 ;
      RECT  8.55 2.62 8.78 3.245 ;
      RECT  8.44 3.245 8.78 3.475 ;
      RECT  10.08 2.1 10.745 2.38 ;
      RECT  10.515 2.38 10.745 2.675 ;
      RECT  14.445 1.65 14.675 2.39 ;
      RECT  14.445 2.39 16.41 2.62 ;
      RECT  14.445 2.62 14.675 3.525 ;
      RECT  7.98 2.335 8.32 2.675 ;
      RECT  7.98 2.675 8.21 3.495 ;
      RECT  4.92 1.29 5.98 1.295 ;
      RECT  4.92 1.295 5.985 1.3 ;
      RECT  4.92 1.3 5.99 1.305 ;
      RECT  4.92 1.305 5.995 1.31 ;
      RECT  4.92 1.31 6.0 1.315 ;
      RECT  4.92 1.315 6.005 1.32 ;
      RECT  4.92 1.32 6.01 1.325 ;
      RECT  4.92 1.325 6.015 1.33 ;
      RECT  4.92 1.33 6.02 1.335 ;
      RECT  4.92 1.335 6.025 1.34 ;
      RECT  4.92 1.34 6.03 1.345 ;
      RECT  4.92 1.345 6.035 1.35 ;
      RECT  4.92 1.35 6.04 1.355 ;
      RECT  4.92 1.355 6.045 1.36 ;
      RECT  4.92 1.36 6.05 1.365 ;
      RECT  4.92 1.365 6.055 1.37 ;
      RECT  4.92 1.37 6.06 1.375 ;
      RECT  4.92 1.375 6.065 1.38 ;
      RECT  4.92 1.38 6.07 1.385 ;
      RECT  4.92 1.385 6.075 1.39 ;
      RECT  4.92 1.39 6.08 1.395 ;
      RECT  4.92 1.395 6.085 1.4 ;
      RECT  4.92 1.4 6.09 1.405 ;
      RECT  4.92 1.405 6.095 1.41 ;
      RECT  4.92 1.41 6.1 1.415 ;
      RECT  4.92 1.415 6.105 1.42 ;
      RECT  4.92 1.42 6.11 1.425 ;
      RECT  4.92 1.425 6.115 1.43 ;
      RECT  4.92 1.43 6.12 1.435 ;
      RECT  4.92 1.435 6.125 1.44 ;
      RECT  4.92 1.44 6.13 1.445 ;
      RECT  4.92 1.445 6.135 1.45 ;
      RECT  4.92 1.45 6.14 1.455 ;
      RECT  4.92 1.455 6.145 1.46 ;
      RECT  4.92 1.46 6.15 1.465 ;
      RECT  4.92 1.465 6.155 1.47 ;
      RECT  4.92 1.47 6.16 1.475 ;
      RECT  4.92 1.475 6.165 1.48 ;
      RECT  4.92 1.48 6.17 1.485 ;
      RECT  4.92 1.485 6.175 1.49 ;
      RECT  4.92 1.49 6.18 1.52 ;
      RECT  5.875 1.52 6.18 1.525 ;
      RECT  4.92 1.52 5.15 1.565 ;
      RECT  5.88 1.525 6.18 1.53 ;
      RECT  5.885 1.53 6.18 1.535 ;
      RECT  5.89 1.535 6.18 1.54 ;
      RECT  5.895 1.54 6.18 1.545 ;
      RECT  5.9 1.545 6.18 1.55 ;
      RECT  5.905 1.55 6.18 1.555 ;
      RECT  5.91 1.555 6.18 1.56 ;
      RECT  5.915 1.56 6.18 1.565 ;
      RECT  2.42 1.565 5.15 1.795 ;
      RECT  5.92 1.565 6.18 1.57 ;
      RECT  5.925 1.57 6.18 1.575 ;
      RECT  5.93 1.575 6.18 1.58 ;
      RECT  5.935 1.58 6.18 1.585 ;
      RECT  5.94 1.585 6.18 1.59 ;
      RECT  5.945 1.59 6.18 1.595 ;
      RECT  5.95 1.595 6.18 3.495 ;
      RECT  2.685 1.795 2.915 3.035 ;
      RECT  2.42 3.035 2.915 3.265 ;
      RECT  5.95 3.495 8.21 3.725 ;
      RECT  3.245 3.955 5.0 4.185 ;
      RECT  3.245 4.185 3.475 4.365 ;
      RECT  4.34 0.83 6.67 1.005 ;
      RECT  0.995 1.005 6.67 1.06 ;
      RECT  6.2 1.06 6.67 1.12 ;
      RECT  0.995 1.06 4.62 1.235 ;
      RECT  6.44 1.12 6.67 2.1 ;
      RECT  1.005 1.235 1.235 3.955 ;
      RECT  6.44 2.1 7.0 2.38 ;
      RECT  0.18 3.955 2.355 4.185 ;
      RECT  2.125 4.185 2.355 4.365 ;
      RECT  2.125 4.365 3.475 4.595 ;
      RECT  0.5 4.415 1.795 4.645 ;
      RECT  0.5 4.645 0.73 5.0 ;
      RECT  1.565 4.645 1.795 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  1.565 5.0 2.97 5.23 ;
      RECT  7.22 4.415 11.315 4.645 ;
      RECT  11.085 4.645 11.315 4.675 ;
      RECT  7.22 4.645 7.45 5.0 ;
      RECT  11.085 4.675 14.06 4.905 ;
      RECT  13.83 4.905 14.06 5.0 ;
      RECT  4.87 5.0 7.45 5.23 ;
      RECT  13.83 5.0 14.17 5.23 ;
      LAYER METAL2 ;
      RECT  6.44 2.1 10.64 2.38 ;
      LAYER VIA12 ;
      RECT  6.59 2.11 6.85 2.37 ;
      RECT  10.23 2.11 10.49 2.37 ;
  END
END MDN_ADDF_P1_2
#-----------------------------------------------------------------------
#      Cell        : MDN_ADDF_P1_4
#      Description : Full adder
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ADDF_P1_4
  CLASS CORE ;
  FOREIGN MDN_ADDF_P1_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 24.64 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 3.49 ;
      RECT  1.54 3.49 4.06 3.72 ;
      RECT  3.78 2.125 4.06 3.49 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  20.34 1.565 24.46 1.795 ;
      RECT  22.285 1.795 22.515 3.245 ;
      RECT  20.34 3.245 24.46 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.86 1.565 19.98 1.795 ;
      RECT  17.805 1.795 18.035 3.245 ;
      RECT  15.86 3.245 19.98 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.81 5.74 ;
      RECT  21.165 4.87 21.395 5.46 ;
      RECT  20.72 5.46 21.395 5.74 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.685 5.46 19.155 5.74 ;
      RECT  18.925 4.87 19.155 5.46 ;
      RECT  9.965 4.93 10.195 5.46 ;
      RECT  9.965 5.46 12.88 5.74 ;
      RECT  12.15 5.135 12.49 5.46 ;
      RECT  7.725 4.93 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.805 4.48 4.3 4.71 ;
      RECT  3.805 4.71 4.035 5.46 ;
      RECT  3.805 5.46 4.48 5.74 ;
      RECT  1.005 4.945 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 24.64 5.74 ;
      LAYER VIA12 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  24.23 5.47 24.49 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  18.07 5.47 18.33 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 -0.14 24.81 0.14 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.52 ;
      RECT  9.405 -0.14 10.08 0.14 ;
      RECT  9.405 0.14 9.635 0.89 ;
      RECT  9.14 0.89 9.635 1.12 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 24.64 0.14 ;
      LAYER VIA12 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  12.665 0.37 15.29 0.6 ;
      RECT  12.665 0.6 12.895 0.75 ;
      RECT  9.965 0.75 12.895 0.98 ;
      RECT  9.965 0.98 10.195 1.35 ;
      RECT  5.99 0.37 7.185 0.6 ;
      RECT  6.955 0.6 7.185 1.29 ;
      RECT  6.955 1.29 8.985 1.295 ;
      RECT  6.955 1.295 8.99 1.3 ;
      RECT  6.955 1.3 8.995 1.305 ;
      RECT  6.955 1.305 9.0 1.31 ;
      RECT  6.955 1.31 9.005 1.315 ;
      RECT  6.955 1.315 9.01 1.32 ;
      RECT  6.955 1.32 9.015 1.325 ;
      RECT  6.955 1.325 9.02 1.33 ;
      RECT  6.955 1.33 9.025 1.335 ;
      RECT  6.955 1.335 9.03 1.34 ;
      RECT  6.955 1.34 9.035 1.345 ;
      RECT  6.955 1.345 9.04 1.35 ;
      RECT  6.955 1.35 10.195 1.52 ;
      RECT  8.88 1.52 10.195 1.525 ;
      RECT  7.165 1.52 7.395 3.03 ;
      RECT  8.885 1.525 10.195 1.53 ;
      RECT  8.89 1.53 10.195 1.535 ;
      RECT  8.895 1.535 10.195 1.54 ;
      RECT  8.9 1.54 10.195 1.545 ;
      RECT  8.905 1.545 10.195 1.55 ;
      RECT  8.91 1.55 10.195 1.555 ;
      RECT  8.915 1.555 10.195 1.56 ;
      RECT  8.92 1.56 10.195 1.565 ;
      RECT  8.925 1.565 10.195 1.57 ;
      RECT  8.93 1.57 10.195 1.575 ;
      RECT  8.935 1.575 10.195 1.58 ;
      RECT  6.9 3.03 7.395 3.26 ;
      RECT  21.67 0.37 23.13 0.6 ;
      RECT  13.125 0.89 13.96 1.12 ;
      RECT  13.125 1.12 13.355 1.29 ;
      RECT  11.38 1.29 13.355 1.52 ;
      RECT  12.205 1.52 12.435 2.415 ;
      RECT  12.205 2.415 13.05 2.645 ;
      RECT  12.205 2.645 12.435 3.245 ;
      RECT  11.38 3.245 12.435 3.475 ;
      RECT  12.205 3.475 12.435 3.755 ;
      RECT  12.205 3.755 15.455 3.76 ;
      RECT  12.205 3.76 15.5 3.985 ;
      RECT  15.16 3.985 15.5 3.99 ;
      RECT  14.19 1.005 15.5 1.235 ;
      RECT  14.19 1.235 14.42 1.295 ;
      RECT  14.185 1.295 14.42 1.3 ;
      RECT  14.18 1.3 14.42 1.305 ;
      RECT  14.175 1.305 14.42 1.31 ;
      RECT  14.17 1.31 14.42 1.315 ;
      RECT  14.165 1.315 14.42 1.32 ;
      RECT  14.16 1.32 14.42 1.325 ;
      RECT  14.155 1.325 14.42 1.33 ;
      RECT  14.15 1.33 14.42 1.335 ;
      RECT  14.145 1.335 14.42 1.34 ;
      RECT  14.14 1.34 14.42 1.345 ;
      RECT  14.135 1.345 14.42 1.35 ;
      RECT  14.13 1.35 14.42 1.355 ;
      RECT  14.125 1.355 14.42 1.36 ;
      RECT  14.12 1.36 14.42 1.365 ;
      RECT  14.115 1.365 14.42 1.37 ;
      RECT  14.11 1.37 14.42 1.375 ;
      RECT  14.105 1.375 14.42 1.38 ;
      RECT  14.1 1.38 14.42 1.385 ;
      RECT  14.095 1.385 14.42 1.39 ;
      RECT  14.09 1.39 14.415 1.395 ;
      RECT  14.085 1.395 14.41 1.4 ;
      RECT  14.08 1.4 14.405 1.405 ;
      RECT  14.075 1.405 14.4 1.41 ;
      RECT  14.07 1.41 14.395 1.415 ;
      RECT  14.065 1.415 14.39 1.42 ;
      RECT  14.06 1.42 14.385 1.425 ;
      RECT  14.055 1.425 14.38 1.43 ;
      RECT  14.05 1.43 14.375 1.435 ;
      RECT  14.045 1.435 14.37 1.44 ;
      RECT  14.04 1.44 14.365 1.445 ;
      RECT  14.035 1.445 14.36 1.45 ;
      RECT  14.03 1.45 14.355 1.455 ;
      RECT  14.025 1.455 14.35 1.46 ;
      RECT  14.02 1.46 14.345 1.465 ;
      RECT  14.015 1.465 14.34 1.47 ;
      RECT  14.01 1.47 14.335 1.475 ;
      RECT  14.005 1.475 14.33 1.48 ;
      RECT  14.0 1.48 14.325 1.485 ;
      RECT  13.995 1.485 14.32 1.49 ;
      RECT  13.99 1.49 14.315 1.495 ;
      RECT  13.985 1.495 14.31 1.5 ;
      RECT  13.98 1.5 14.305 1.505 ;
      RECT  13.975 1.505 14.3 1.51 ;
      RECT  13.97 1.51 14.295 1.515 ;
      RECT  13.97 1.515 14.29 1.52 ;
      RECT  13.97 1.52 14.285 1.525 ;
      RECT  13.97 1.525 14.28 1.53 ;
      RECT  13.97 1.53 14.275 1.535 ;
      RECT  13.97 1.535 14.27 1.54 ;
      RECT  13.97 1.54 14.265 1.545 ;
      RECT  13.97 1.545 14.26 1.55 ;
      RECT  13.97 1.55 14.255 1.555 ;
      RECT  13.97 1.555 14.25 1.56 ;
      RECT  13.97 1.56 14.245 1.565 ;
      RECT  13.97 1.565 14.24 1.57 ;
      RECT  13.97 1.57 14.235 1.575 ;
      RECT  13.97 1.575 14.23 1.58 ;
      RECT  13.97 1.58 14.225 1.585 ;
      RECT  13.97 1.585 14.22 1.59 ;
      RECT  13.97 1.59 14.215 1.595 ;
      RECT  13.97 1.595 14.21 1.6 ;
      RECT  13.97 1.6 14.205 1.605 ;
      RECT  13.97 1.605 14.2 1.75 ;
      RECT  12.92 1.75 14.2 1.98 ;
      RECT  13.325 1.98 13.555 3.245 ;
      RECT  12.92 3.245 13.96 3.475 ;
      RECT  10.68 1.565 11.15 1.795 ;
      RECT  10.92 1.795 11.15 2.41 ;
      RECT  10.92 2.41 11.93 2.64 ;
      RECT  10.92 2.64 11.15 3.245 ;
      RECT  9.14 3.245 11.15 3.475 ;
      RECT  5.43 1.75 5.77 1.98 ;
      RECT  5.485 1.98 5.715 3.95 ;
      RECT  5.485 3.95 11.875 4.18 ;
      RECT  11.645 4.18 11.875 4.215 ;
      RECT  11.645 4.215 14.675 4.365 ;
      RECT  11.645 4.365 21.9 4.445 ;
      RECT  14.445 4.445 21.9 4.595 ;
      RECT  20.55 4.595 20.78 5.0 ;
      RECT  21.67 4.595 21.9 5.0 ;
      RECT  20.55 5.0 20.89 5.23 ;
      RECT  21.67 5.0 22.01 5.23 ;
      RECT  8.44 1.75 8.78 1.98 ;
      RECT  8.55 1.98 8.78 2.4 ;
      RECT  8.55 2.4 9.69 2.63 ;
      RECT  8.55 2.63 8.78 3.245 ;
      RECT  8.44 3.245 8.78 3.475 ;
      RECT  10.08 2.1 10.69 2.38 ;
      RECT  10.46 2.38 10.69 2.685 ;
      RECT  14.445 1.695 14.675 2.395 ;
      RECT  14.445 2.395 17.53 2.625 ;
      RECT  14.445 2.625 14.675 3.245 ;
      RECT  14.39 3.245 14.73 3.475 ;
      RECT  8.09 2.355 8.32 2.465 ;
      RECT  7.725 2.465 8.32 2.695 ;
      RECT  7.725 2.695 7.955 3.49 ;
      RECT  4.925 1.29 5.975 1.295 ;
      RECT  4.925 1.295 5.98 1.3 ;
      RECT  4.925 1.3 5.985 1.305 ;
      RECT  4.925 1.305 5.99 1.31 ;
      RECT  4.925 1.31 5.995 1.315 ;
      RECT  4.925 1.315 6.0 1.32 ;
      RECT  4.925 1.32 6.005 1.325 ;
      RECT  4.925 1.325 6.01 1.33 ;
      RECT  4.925 1.33 6.015 1.335 ;
      RECT  4.925 1.335 6.02 1.34 ;
      RECT  4.925 1.34 6.025 1.345 ;
      RECT  4.925 1.345 6.03 1.35 ;
      RECT  4.925 1.35 6.035 1.355 ;
      RECT  4.925 1.355 6.04 1.36 ;
      RECT  4.925 1.36 6.045 1.365 ;
      RECT  4.925 1.365 6.05 1.37 ;
      RECT  4.925 1.37 6.055 1.375 ;
      RECT  4.925 1.375 6.06 1.38 ;
      RECT  4.925 1.38 6.065 1.385 ;
      RECT  4.925 1.385 6.07 1.39 ;
      RECT  4.925 1.39 6.075 1.395 ;
      RECT  4.925 1.395 6.08 1.4 ;
      RECT  4.925 1.4 6.085 1.405 ;
      RECT  4.925 1.405 6.09 1.41 ;
      RECT  4.925 1.41 6.095 1.415 ;
      RECT  4.925 1.415 6.1 1.42 ;
      RECT  4.925 1.42 6.105 1.425 ;
      RECT  4.925 1.425 6.11 1.43 ;
      RECT  4.925 1.43 6.115 1.435 ;
      RECT  4.925 1.435 6.12 1.44 ;
      RECT  4.925 1.44 6.125 1.445 ;
      RECT  4.925 1.445 6.13 1.45 ;
      RECT  4.925 1.45 6.135 1.455 ;
      RECT  4.925 1.455 6.14 1.46 ;
      RECT  4.925 1.46 6.145 1.465 ;
      RECT  4.925 1.465 6.15 1.47 ;
      RECT  4.925 1.47 6.155 1.475 ;
      RECT  4.925 1.475 6.16 1.48 ;
      RECT  4.925 1.48 6.165 1.485 ;
      RECT  4.925 1.485 6.17 1.49 ;
      RECT  4.925 1.49 6.175 1.495 ;
      RECT  4.925 1.495 6.18 1.5 ;
      RECT  4.925 1.5 6.185 1.505 ;
      RECT  4.925 1.505 6.19 1.51 ;
      RECT  4.925 1.51 6.195 1.515 ;
      RECT  4.925 1.515 6.2 1.52 ;
      RECT  5.87 1.52 6.205 1.525 ;
      RECT  4.925 1.52 5.155 1.565 ;
      RECT  5.875 1.525 6.21 1.53 ;
      RECT  5.88 1.53 6.215 1.535 ;
      RECT  5.885 1.535 6.22 1.54 ;
      RECT  5.89 1.54 6.225 1.545 ;
      RECT  5.895 1.545 6.23 1.55 ;
      RECT  5.9 1.55 6.23 1.555 ;
      RECT  5.905 1.555 6.23 1.56 ;
      RECT  5.91 1.56 6.23 1.565 ;
      RECT  2.42 1.565 5.155 1.795 ;
      RECT  5.915 1.565 6.23 1.57 ;
      RECT  5.92 1.57 6.23 1.575 ;
      RECT  5.925 1.575 6.23 1.58 ;
      RECT  5.93 1.58 6.23 1.585 ;
      RECT  5.935 1.585 6.23 1.59 ;
      RECT  5.94 1.59 6.23 1.595 ;
      RECT  5.945 1.595 6.23 1.6 ;
      RECT  5.95 1.6 6.23 1.605 ;
      RECT  5.955 1.605 6.23 1.61 ;
      RECT  5.96 1.61 6.23 1.615 ;
      RECT  5.965 1.615 6.23 1.62 ;
      RECT  5.97 1.62 6.23 1.625 ;
      RECT  5.975 1.625 6.23 1.63 ;
      RECT  5.98 1.63 6.23 1.635 ;
      RECT  5.985 1.635 6.23 1.64 ;
      RECT  5.99 1.64 6.23 1.645 ;
      RECT  5.995 1.645 6.23 1.65 ;
      RECT  6.0 1.65 6.23 3.49 ;
      RECT  2.685 1.795 2.915 3.03 ;
      RECT  2.42 3.03 2.915 3.26 ;
      RECT  6.0 3.49 7.955 3.72 ;
      RECT  22.79 2.405 24.25 2.635 ;
      RECT  18.31 2.41 19.77 2.64 ;
      RECT  3.245 4.02 5.0 4.25 ;
      RECT  3.245 4.25 3.475 4.365 ;
      RECT  4.365 0.83 6.69 1.005 ;
      RECT  1.005 1.005 6.69 1.06 ;
      RECT  6.2 1.06 6.69 1.12 ;
      RECT  1.005 1.06 4.595 1.235 ;
      RECT  6.46 1.12 6.69 2.1 ;
      RECT  1.005 1.235 1.235 3.95 ;
      RECT  6.46 2.1 6.84 2.38 ;
      RECT  0.18 3.95 2.355 4.18 ;
      RECT  2.125 4.18 2.355 4.365 ;
      RECT  2.125 4.365 3.475 4.595 ;
      RECT  7.22 4.41 11.315 4.64 ;
      RECT  11.085 4.64 11.315 4.675 ;
      RECT  7.22 4.64 7.45 5.0 ;
      RECT  11.085 4.675 14.06 4.905 ;
      RECT  13.83 4.905 14.06 5.0 ;
      RECT  4.87 5.0 7.45 5.23 ;
      RECT  13.83 5.0 14.17 5.23 ;
      RECT  0.5 4.485 1.795 4.715 ;
      RECT  0.5 4.715 0.75 5.0 ;
      RECT  1.49 4.715 1.795 5.0 ;
      RECT  0.39 5.0 0.75 5.23 ;
      RECT  1.49 5.0 2.97 5.23 ;
      RECT  17.19 5.0 18.65 5.23 ;
      LAYER METAL2 ;
      RECT  6.46 2.1 10.69 2.38 ;
      LAYER VIA12 ;
      RECT  6.52 2.11 6.78 2.37 ;
      RECT  10.37 2.11 10.63 2.37 ;
  END
END MDN_ADDF_P1_4
#-----------------------------------------------------------------------
#      Cell        : MDN_ADDH_1
#      Description : Half adder
#      Equation    : S=A^B:CO=A&B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ADDH_1
  CLASS CORE ;
  FOREIGN MDN_ADDH_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.565 2.115 2.9 2.125 ;
      RECT  1.54 2.125 2.94 2.345 ;
      RECT  1.54 2.345 1.82 2.915 ;
      RECT  2.66 2.345 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 7.395 1.795 ;
      RECT  7.165 1.795 7.395 3.245 ;
      RECT  6.9 3.245 7.395 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.285 1.565 8.78 1.795 ;
      RECT  8.285 1.795 8.515 3.245 ;
      RECT  8.285 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 4.365 6.54 4.595 ;
      RECT  6.045 4.595 6.275 5.46 ;
      RECT  6.045 5.46 7.955 5.74 ;
      RECT  7.725 4.905 7.955 5.46 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.905 1.235 5.46 ;
      RECT  0.56 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  4.48 -0.14 5.155 0.14 ;
      RECT  4.925 0.14 5.155 1.005 ;
      RECT  4.66 1.005 5.155 1.235 ;
      RECT  1.565 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.695 ;
      RECT  1.565 0.14 1.795 1.005 ;
      RECT  1.565 1.005 2.06 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  0.18 1.005 1.23 1.235 ;
      RECT  1.0 1.235 1.23 1.565 ;
      RECT  1.0 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 2.125 ;
      RECT  1.0 1.795 1.23 3.805 ;
      RECT  3.245 2.125 6.05 2.355 ;
      RECT  5.82 2.355 6.05 2.69 ;
      RECT  0.18 3.805 2.06 4.035 ;
      RECT  2.42 1.005 4.035 1.235 ;
      RECT  3.805 1.235 4.035 1.565 ;
      RECT  3.805 1.565 5.77 1.795 ;
      RECT  6.2 1.565 6.595 1.795 ;
      RECT  6.365 1.795 6.595 3.245 ;
      RECT  5.43 3.245 6.595 3.475 ;
      RECT  6.365 3.475 6.595 3.805 ;
      RECT  6.365 3.805 7.395 4.035 ;
      RECT  7.165 4.035 7.395 4.365 ;
      RECT  7.165 4.365 8.45 4.595 ;
      RECT  8.22 4.595 8.45 5.0 ;
      RECT  8.22 5.0 8.57 5.23 ;
      RECT  2.42 3.805 4.595 4.035 ;
      RECT  4.365 4.035 4.595 4.365 ;
      RECT  4.365 4.365 5.0 4.595 ;
      RECT  0.5 4.365 4.035 4.595 ;
      RECT  0.5 4.595 0.73 5.0 ;
      RECT  3.805 4.595 4.035 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  3.805 5.0 5.21 5.23 ;
  END
END MDN_ADDH_1
#-----------------------------------------------------------------------
#      Cell        : MDN_ADDH_2
#      Description : Half adder
#      Equation    : S=A^B:CO=A&B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ADDH_2
  CLASS CORE ;
  FOREIGN MDN_ADDH_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.545 2.115 2.92 2.125 ;
      RECT  1.54 2.125 2.94 2.345 ;
      RECT  1.54 2.345 1.82 2.915 ;
      RECT  2.66 2.345 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 8.78 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  6.875 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.135 1.565 11.02 1.795 ;
      RECT  9.965 1.795 10.195 3.245 ;
      RECT  9.14 3.245 11.02 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  6.2 4.365 6.835 4.595 ;
      RECT  6.605 4.595 6.835 5.46 ;
      RECT  6.55 5.46 7.955 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  3.245 4.905 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.905 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  1.565 -0.14 4.65 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  1.565 0.14 1.795 1.005 ;
      RECT  4.365 0.14 4.595 1.005 ;
      RECT  1.565 1.005 2.06 1.235 ;
      RECT  4.365 1.005 5.0 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 8.57 0.6 ;
      RECT  8.23 0.6 8.46 1.005 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  7.22 0.6 7.45 1.005 ;
      RECT  7.22 1.005 8.46 1.125 ;
      RECT  7.225 1.125 8.46 1.235 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 1.565 ;
      RECT  1.005 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 2.125 ;
      RECT  1.005 1.795 1.235 3.805 ;
      RECT  3.245 2.125 6.05 2.355 ;
      RECT  5.82 2.355 6.05 2.69 ;
      RECT  0.18 3.805 2.06 4.035 ;
      RECT  2.42 1.005 4.035 1.235 ;
      RECT  3.805 1.235 4.035 1.565 ;
      RECT  3.805 1.565 5.77 1.795 ;
      RECT  6.2 1.565 6.595 1.795 ;
      RECT  6.365 1.795 6.595 3.245 ;
      RECT  5.43 3.245 6.595 3.475 ;
      RECT  6.365 3.475 6.595 3.805 ;
      RECT  6.365 3.805 7.395 4.035 ;
      RECT  7.165 4.035 7.395 4.365 ;
      RECT  7.165 4.365 10.7 4.595 ;
      RECT  9.46 4.595 9.69 5.0 ;
      RECT  10.47 4.595 10.7 5.0 ;
      RECT  9.35 5.0 9.69 5.23 ;
      RECT  10.47 5.0 10.81 5.23 ;
      RECT  2.42 3.805 4.595 4.035 ;
      RECT  4.365 4.035 4.595 4.365 ;
      RECT  4.365 4.365 5.0 4.595 ;
      RECT  0.445 4.355 4.035 4.365 ;
      RECT  0.42 4.365 4.035 4.585 ;
      RECT  0.42 4.585 0.7 5.0 ;
      RECT  3.805 4.585 4.035 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  3.805 5.0 5.21 5.23 ;
  END
END MDN_ADDH_2
#-----------------------------------------------------------------------
#      Cell        : MDN_ADDH_4
#      Description : Half adder
#      Equation    : S=A^B:CO=A&B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ADDH_4
  CLASS CORE ;
  FOREIGN MDN_ADDH_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.545 2.115 2.92 2.125 ;
      RECT  1.54 2.125 2.94 2.345 ;
      RECT  1.54 2.345 1.82 2.915 ;
      RECT  2.66 2.345 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 11.02 1.795 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  6.875 3.245 11.02 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.38 1.565 15.5 1.795 ;
      RECT  14.445 1.795 14.675 3.245 ;
      RECT  11.355 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.93 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.93 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.965 4.93 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  6.045 4.365 6.54 4.595 ;
      RECT  6.045 4.595 6.275 5.46 ;
      RECT  6.045 5.46 7.955 5.74 ;
      RECT  7.725 4.93 7.955 5.46 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.695 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  12.205 0.14 12.435 0.695 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  4.48 -0.14 5.155 0.14 ;
      RECT  4.925 0.14 5.155 1.005 ;
      RECT  4.66 1.005 5.155 1.235 ;
      RECT  1.565 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.695 ;
      RECT  1.565 0.14 1.795 1.005 ;
      RECT  1.565 1.005 2.06 1.235 ;
      RECT  -0.17 -0.14 0.65 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  8.22 0.37 9.69 0.6 ;
      RECT  14.94 0.37 15.28 0.6 ;
      RECT  14.94 0.6 15.17 1.005 ;
      RECT  12.7 0.37 13.04 0.375 ;
      RECT  12.7 0.375 14.17 0.605 ;
      RECT  13.83 0.37 14.17 0.375 ;
      RECT  12.7 0.605 12.93 1.005 ;
      RECT  13.94 0.605 14.17 1.005 ;
      RECT  10.525 0.37 11.955 0.6 ;
      RECT  10.525 0.6 10.755 1.005 ;
      RECT  11.725 0.6 11.955 1.005 ;
      RECT  6.365 1.005 10.755 1.235 ;
      RECT  11.725 1.005 12.93 1.235 ;
      RECT  13.94 1.005 15.17 1.235 ;
      RECT  6.365 1.235 6.595 1.565 ;
      RECT  6.2 1.565 6.595 1.795 ;
      RECT  6.365 1.795 6.595 3.245 ;
      RECT  5.43 3.245 6.595 3.475 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 1.565 ;
      RECT  1.005 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 2.125 ;
      RECT  1.005 1.795 1.235 3.805 ;
      RECT  3.245 2.125 6.05 2.355 ;
      RECT  5.82 2.355 6.05 2.69 ;
      RECT  0.18 3.805 2.06 4.035 ;
      RECT  2.42 1.005 4.035 1.235 ;
      RECT  3.805 1.235 4.035 1.565 ;
      RECT  3.805 1.565 5.77 1.795 ;
      RECT  7.165 2.335 7.395 2.685 ;
      RECT  7.165 2.685 8.515 2.915 ;
      RECT  8.285 2.335 8.515 2.685 ;
      RECT  9.405 2.35 9.635 2.685 ;
      RECT  9.405 2.685 10.755 2.915 ;
      RECT  10.525 2.35 10.755 2.685 ;
      RECT  2.42 3.805 4.595 4.035 ;
      RECT  4.365 4.035 4.595 4.365 ;
      RECT  4.365 4.365 5.0 4.595 ;
      RECT  0.5 4.365 4.035 4.595 ;
      RECT  0.5 4.595 0.73 5.0 ;
      RECT  3.805 4.595 4.035 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  3.805 5.0 5.21 5.23 ;
  END
END MDN_ADDH_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AN2_1
#      Description : 2-Input AND
#      Equation    : X=A1&A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN2_1
  CLASS CORE ;
  FOREIGN MDN_AN2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.695 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 3.805 ;
      RECT  2.42 3.805 3.475 4.035 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  1.565 3.245 2.915 3.475 ;
      RECT  1.565 3.475 1.795 3.805 ;
      RECT  0.18 3.805 1.795 4.035 ;
  END
END MDN_AN2_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AN2_12
#      Description : 2-Input AND
#      Equation    : X=A1&A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN2_12
  CLASS CORE ;
  FOREIGN MDN_AN2_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.685 ;
      RECT  3.78 2.685 6.3 2.915 ;
      RECT  4.9 2.125 5.18 2.685 ;
      RECT  6.02 2.125 6.3 2.685 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.93 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.93 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  12.205 4.93 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 4.93 14.675 5.46 ;
      RECT  9.965 4.93 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.67 4.985 8.01 5.46 ;
      RECT  7.28 5.46 8.4 5.74 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.695 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.695 ;
      RECT  12.205 -0.14 14.675 0.14 ;
      RECT  12.205 0.14 12.435 0.695 ;
      RECT  14.445 0.14 14.675 0.695 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.67 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 2.76 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.955 0.92 8.04 1.32 ;
      RECT  7.64 1.32 8.04 1.54 ;
      RECT  7.64 1.54 19.925 1.94 ;
      RECT  17.715 1.94 18.115 3.1 ;
      RECT  7.725 3.1 19.925 3.105 ;
      RECT  7.64 3.105 19.925 3.5 ;
      RECT  7.64 3.5 8.04 4.28 ;
      RECT  6.96 4.28 8.04 4.31 ;
      RECT  6.955 4.31 8.04 4.65 ;
      RECT  6.96 4.65 8.04 4.68 ;
    END
    ANTENNADIFFAREA 18.144 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  19.42 0.37 19.77 0.6 ;
      RECT  19.42 0.6 19.65 1.005 ;
      RECT  17.19 0.37 18.65 0.6 ;
      RECT  18.42 0.6 18.65 1.005 ;
      RECT  18.42 1.005 19.65 1.235 ;
      RECT  0.95 0.445 5.77 0.675 ;
      RECT  3.91 1.005 6.275 1.235 ;
      RECT  6.045 1.235 6.275 1.565 ;
      RECT  6.045 1.565 7.395 1.795 ;
      RECT  7.165 1.795 7.395 2.405 ;
      RECT  7.165 2.405 17.485 2.635 ;
      RECT  7.165 2.635 7.395 3.805 ;
      RECT  6.045 3.805 7.395 4.035 ;
      RECT  6.045 4.035 6.275 4.365 ;
      RECT  0.14 4.365 6.275 4.595 ;
  END
END MDN_AN2_12
#-----------------------------------------------------------------------
#      Cell        : MDN_AN2_2
#      Description : 2-Input AND
#      Equation    : X=A1&A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN2_2
  CLASS CORE ;
  FOREIGN MDN_AN2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.645 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 0.945 ;
      RECT  0.18 0.945 0.675 1.175 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 4.3 1.795 ;
      RECT  3.245 1.795 3.475 3.245 ;
      RECT  2.42 3.245 4.3 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.74 0.37 4.08 0.6 ;
      RECT  3.74 0.6 3.97 1.005 ;
      RECT  2.63 0.37 2.97 0.6 ;
      RECT  2.74 0.6 2.97 1.005 ;
      RECT  1.005 1.005 3.97 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 2.06 4.595 ;
  END
END MDN_AN2_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AN2_3
#      Description : 2-Input AND
#      Equation    : X=A1&A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN2_3
  CLASS CORE ;
  FOREIGN MDN_AN2_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  3.245 5.46 5.715 5.74 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.58 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.58 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.125 1.005 2.9 1.235 ;
      RECT  2.67 1.235 2.9 1.565 ;
      RECT  2.67 1.565 5.0 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  2.67 3.245 5.0 3.475 ;
      RECT  2.67 3.475 2.9 4.365 ;
      RECT  2.42 4.365 2.9 4.595 ;
    END
    ANTENNADIFFAREA 4.536 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.67 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 2.405 ;
      RECT  2.125 2.405 4.09 2.635 ;
      RECT  2.125 2.635 2.355 3.805 ;
      RECT  1.565 3.805 2.355 4.035 ;
      RECT  1.565 4.035 1.795 4.365 ;
      RECT  0.18 4.365 1.795 4.595 ;
      RECT  3.75 5.0 5.21 5.23 ;
  END
END MDN_AN2_3
#-----------------------------------------------------------------------
#      Cell        : MDN_AN2_4
#      Description : 2-Input AND
#      Equation    : X=A1&A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN2_4
  CLASS CORE ;
  FOREIGN MDN_AN2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.585 ;
      RECT  5.485 0.14 5.715 0.585 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  3.245 1.565 6.54 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  3.805 3.245 6.54 3.475 ;
      RECT  3.805 3.475 4.035 3.805 ;
      RECT  2.42 3.805 4.035 4.035 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.985 0.37 6.33 0.6 ;
      RECT  5.985 0.6 6.215 1.005 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  4.98 1.005 6.215 1.235 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 2.38 ;
      RECT  2.685 2.38 5.12 2.61 ;
      RECT  2.685 2.61 2.915 3.245 ;
      RECT  1.565 3.245 2.915 3.475 ;
      RECT  1.565 3.475 1.795 3.805 ;
      RECT  0.18 3.805 1.795 4.035 ;
  END
END MDN_AN2_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AN2_6
#      Description : 2-Input AND
#      Equation    : X=A1&A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN2_6
  CLASS CORE ;
  FOREIGN MDN_AN2_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.67 2.115 3.995 2.125 ;
      RECT  2.66 2.125 4.06 2.345 ;
      RECT  2.66 2.345 2.94 2.915 ;
      RECT  3.78 2.345 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.43 2.115 1.755 2.125 ;
      RECT  0.42 2.125 1.82 2.345 ;
      RECT  0.42 2.345 0.7 2.915 ;
      RECT  1.54 2.345 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.93 7.955 5.46 ;
      RECT  7.725 5.46 11.37 5.74 ;
      RECT  9.965 4.93 10.195 5.46 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.58 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.005 5.155 1.235 ;
      RECT  4.925 1.235 5.155 1.565 ;
      RECT  4.925 1.565 11.02 1.795 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  4.925 3.245 11.02 3.475 ;
      RECT  4.925 3.475 5.155 4.365 ;
      RECT  4.66 4.365 5.155 4.595 ;
    END
    ANTENNADIFFAREA 9.072 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.14 1.005 4.3 1.235 ;
      RECT  3.19 1.565 4.595 1.795 ;
      RECT  4.365 1.795 4.595 2.38 ;
      RECT  4.365 2.38 8.475 2.61 ;
      RECT  4.365 2.61 4.595 3.805 ;
      RECT  3.805 3.805 4.595 4.035 ;
      RECT  3.805 4.035 4.035 4.365 ;
      RECT  0.14 4.365 4.035 4.595 ;
      RECT  9.35 2.38 10.81 2.61 ;
      RECT  8.23 5.0 9.69 5.23 ;
  END
END MDN_AN2_6
#-----------------------------------------------------------------------
#      Cell        : MDN_AN2_8
#      Description : 2-Input AND
#      Equation    : X=A1&A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN2_8
  CLASS CORE ;
  FOREIGN MDN_AN2_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.695 ;
      RECT  2.66 2.695 4.06 2.915 ;
      RECT  3.78 2.125 4.06 2.695 ;
      RECT  2.685 2.915 3.9 2.925 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.445 2.115 1.815 2.125 ;
      RECT  0.42 2.125 1.82 2.345 ;
      RECT  0.42 2.345 0.7 2.915 ;
      RECT  1.54 2.345 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.93 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  7.725 4.93 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 4.93 10.195 5.46 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  3.245 5.46 5.715 5.74 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.56 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.585 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.585 ;
      RECT  7.725 0.14 7.955 0.585 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.585 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.005 5.16 1.235 ;
      RECT  4.92 1.235 5.16 1.495 ;
      RECT  4.92 1.495 13.205 1.865 ;
      RECT  12.14 1.865 12.505 3.175 ;
      RECT  4.92 3.175 13.205 3.545 ;
      RECT  4.92 3.545 5.16 3.805 ;
      RECT  4.66 3.805 5.16 4.035 ;
    END
    ANTENNADIFFAREA 12.096 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 0.915 ;
      RECT  11.59 0.37 11.93 0.6 ;
      RECT  11.7 0.6 11.93 0.915 ;
      RECT  11.7 0.915 12.94 1.145 ;
      RECT  1.83 0.445 3.53 0.675 ;
      RECT  1.83 0.675 2.06 1.005 ;
      RECT  0.18 1.005 2.06 1.235 ;
      RECT  2.42 1.005 4.035 1.235 ;
      RECT  3.805 1.235 4.035 1.565 ;
      RECT  3.805 1.565 4.615 1.795 ;
      RECT  4.345 1.795 4.615 2.685 ;
      RECT  4.345 2.685 11.675 2.915 ;
      RECT  4.925 2.35 5.155 2.685 ;
      RECT  6.045 2.35 6.275 2.685 ;
      RECT  7.165 2.35 7.395 2.685 ;
      RECT  8.285 2.35 8.515 2.685 ;
      RECT  9.405 2.35 9.635 2.685 ;
      RECT  10.525 2.35 10.755 2.685 ;
      RECT  11.445 2.35 11.675 2.685 ;
      RECT  4.345 2.915 4.615 3.245 ;
      RECT  3.805 3.245 4.615 3.475 ;
      RECT  3.805 3.475 4.035 3.805 ;
      RECT  0.18 3.805 4.035 4.035 ;
  END
END MDN_AN2_8
#-----------------------------------------------------------------------
#      Cell        : MDN_AN3_1
#      Description : 3-Input AND
#      Equation    : X=A1&A2&A3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN3_1
  CLASS CORE ;
  FOREIGN MDN_AN3_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  1.005 5.46 3.475 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  2.07 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 1.23 1.235 ;
      RECT  1.0 1.235 1.23 1.565 ;
      RECT  1.0 1.565 2.375 1.795 ;
      RECT  2.105 1.795 2.375 4.365 ;
      RECT  0.18 4.365 3.97 4.595 ;
      RECT  3.74 4.595 3.97 5.0 ;
      RECT  3.74 5.0 4.09 5.23 ;
      RECT  1.72 1.005 2.76 1.235 ;
  END
END MDN_AN3_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AN3_2
#      Description : 3-Input AND
#      Equation    : X=A1&A2&A3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN3_2
  CLASS CORE ;
  FOREIGN MDN_AN3_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.905 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.905 1.235 5.46 ;
      RECT  1.005 5.46 3.475 5.74 ;
      RECT  3.245 4.905 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  4.31 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  1.005 -0.14 1.68 0.14 ;
      RECT  1.005 0.14 1.235 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 6.54 1.795 ;
      RECT  5.485 1.795 5.715 3.805 ;
      RECT  4.625 3.805 6.54 4.035 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.98 0.37 6.32 0.6 ;
      RECT  5.98 0.6 6.21 1.005 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  3.245 1.005 6.21 1.235 ;
      RECT  3.245 1.235 3.475 3.805 ;
      RECT  1.715 3.805 4.3 4.035 ;
      RECT  1.715 1.005 2.76 1.235 ;
  END
END MDN_AN3_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AN3_4
#      Description : 3-Input AND
#      Equation    : X=A1&A2&A3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN3_4
  CLASS CORE ;
  FOREIGN MDN_AN3_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.93 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  1.005 5.46 3.475 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  2.07 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.765 1.565 7.37 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  3.785 3.245 7.38 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.985 0.37 7.45 0.6 ;
      RECT  5.985 0.6 6.215 1.005 ;
      RECT  3.74 0.37 5.21 0.6 ;
      RECT  3.74 0.6 3.97 1.005 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  0.43 0.445 2.9 0.675 ;
      RECT  0.43 0.675 0.66 1.005 ;
      RECT  2.67 0.675 2.9 1.005 ;
      RECT  0.18 1.005 0.66 1.235 ;
      RECT  2.67 1.005 3.97 1.235 ;
      RECT  4.98 1.005 6.215 1.235 ;
      RECT  3.245 1.235 3.475 4.365 ;
      RECT  0.18 4.365 3.475 4.595 ;
      RECT  1.72 1.005 2.355 1.235 ;
      RECT  2.125 1.235 2.355 1.565 ;
      RECT  2.125 1.565 2.76 1.795 ;
  END
END MDN_AN3_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AN3_6
#      Description : 3-Input AND
#      Equation    : X=A1&A2&A3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN3_6
  CLASS CORE ;
  FOREIGN MDN_AN3_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.91 2.115 6.235 2.125 ;
      RECT  4.9 2.125 6.3 2.345 ;
      RECT  4.9 2.345 5.18 2.915 ;
      RECT  6.02 2.345 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.67 2.115 3.995 2.125 ;
      RECT  2.66 2.125 4.06 2.345 ;
      RECT  2.66 2.345 2.94 2.915 ;
      RECT  3.78 2.345 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.43 2.115 1.755 2.125 ;
      RECT  0.42 2.125 1.82 2.345 ;
      RECT  0.42 2.345 0.7 2.915 ;
      RECT  1.54 2.345 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.905 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.905 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.93 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.695 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.89 1.005 7.955 1.235 ;
      RECT  7.725 1.235 7.955 1.565 ;
      RECT  7.725 1.565 13.26 1.795 ;
      RECT  11.085 1.795 11.315 3.245 ;
      RECT  7.725 3.245 13.26 3.475 ;
      RECT  7.725 3.475 7.955 4.365 ;
      RECT  6.9 4.365 7.955 4.595 ;
    END
    ANTENNADIFFAREA 9.072 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  12.7 0.37 13.04 0.6 ;
      RECT  12.7 0.6 12.93 1.005 ;
      RECT  10.47 0.37 11.93 0.6 ;
      RECT  11.7 0.6 11.93 1.005 ;
      RECT  11.7 1.005 12.93 1.235 ;
      RECT  3.145 0.445 5.77 0.675 ;
      RECT  0.145 1.005 4.3 1.235 ;
      RECT  4.62 1.005 6.485 1.235 ;
      RECT  6.255 1.235 6.485 1.565 ;
      RECT  6.255 1.565 7.395 1.795 ;
      RECT  7.165 1.795 7.395 2.125 ;
      RECT  7.165 2.125 10.755 2.355 ;
      RECT  8.285 2.355 8.515 2.69 ;
      RECT  9.405 2.355 9.635 2.69 ;
      RECT  10.525 2.355 10.755 2.69 ;
      RECT  7.165 2.355 7.395 3.805 ;
      RECT  6.045 3.805 7.395 4.035 ;
      RECT  6.045 4.035 6.275 4.365 ;
      RECT  0.145 4.365 6.275 4.595 ;
  END
END MDN_AN3_6
#-----------------------------------------------------------------------
#      Cell        : MDN_AN3B_1
#      Description : 3-Input AND (A inverted input)
#      Equation    : X=!A&B1&B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN3B_1
  CLASS CORE ;
  FOREIGN MDN_AN3B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 4.65 5.74 ;
      RECT  1.565 4.365 2.06 4.595 ;
      RECT  1.565 4.595 1.795 5.46 ;
      RECT  1.565 5.46 2.24 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 -0.14 4.65 0.14 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  1.67 1.005 4.3 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  4.07 -0.13 4.33 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.685 1.565 3.53 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  2.42 3.245 2.915 3.475 ;
    END
    ANTENNADIFFAREA 1.992 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.005 0.37 2.97 0.6 ;
      RECT  1.005 0.6 1.235 1.005 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 3.41 ;
  END
END MDN_AN3B_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AN3B_2
#      Description : 3-Input AND (A inverted input)
#      Equation    : X=!A&B1&B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN3B_2
  CLASS CORE ;
  FOREIGN MDN_AN3B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  1.005 5.46 3.475 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.61 ;
      RECT  4.31 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.61 ;
      RECT  0.56 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.005 8.78 1.235 ;
      RECT  5.485 1.235 5.715 3.245 ;
      RECT  4.66 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 4.252 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.83 0.445 3.53 0.675 ;
      RECT  1.83 0.675 2.06 1.005 ;
      RECT  0.145 1.005 2.06 1.235 ;
      RECT  2.42 1.005 4.3 1.235 ;
      RECT  2.42 1.235 2.65 1.575 ;
      RECT  2.125 1.575 2.65 1.805 ;
      RECT  2.125 1.805 2.355 4.365 ;
      RECT  0.18 4.365 4.595 4.595 ;
      RECT  4.365 4.595 4.595 5.0 ;
      RECT  4.365 5.0 6.33 5.23 ;
      RECT  5.43 4.365 8.78 4.595 ;
  END
END MDN_AN3B_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AN3B_3
#      Description : 3-Input AND (A inverted input)
#      Equation    : X=!A&B1&B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN3B_3
  CLASS CORE ;
  FOREIGN MDN_AN3B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.695 ;
      RECT  10.5 2.695 13.02 2.915 ;
      RECT  11.62 2.125 11.9 2.695 ;
      RECT  12.74 2.125 13.02 2.695 ;
      RECT  10.525 2.915 12.955 2.925 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.695 ;
      RECT  3.78 2.695 6.3 2.915 ;
      RECT  4.9 2.125 5.18 2.695 ;
      RECT  6.02 2.125 6.3 2.695 ;
      RECT  3.78 2.915 6.235 2.925 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.43 2.115 2.9 2.125 ;
      RECT  0.42 2.125 2.94 2.345 ;
      RECT  0.42 2.345 0.7 2.915 ;
      RECT  1.54 2.345 1.82 2.915 ;
      RECT  2.66 2.345 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.68 4.365 13.26 4.595 ;
      RECT  12.765 4.595 12.995 5.46 ;
      RECT  12.32 5.46 13.61 5.74 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.695 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.69 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 2.76 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 1.005 13.26 1.235 ;
      RECT  9.965 1.235 10.195 1.565 ;
      RECT  6.9 1.005 7.955 1.235 ;
      RECT  7.725 1.235 7.955 1.565 ;
      RECT  7.725 1.565 10.195 1.795 ;
      RECT  9.965 1.795 10.195 3.245 ;
      RECT  7.725 3.245 10.195 3.475 ;
      RECT  7.725 3.475 7.955 3.805 ;
      RECT  6.9 3.805 7.955 4.035 ;
    END
    ANTENNADIFFAREA 6.378 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 5.77 0.675 ;
      RECT  3.96 1.005 6.275 1.235 ;
      RECT  6.045 1.235 6.275 1.565 ;
      RECT  6.045 1.565 7.395 1.795 ;
      RECT  7.165 1.795 7.395 2.69 ;
      RECT  7.165 2.69 9.635 2.92 ;
      RECT  8.285 2.35 8.515 2.69 ;
      RECT  9.405 2.35 9.635 2.69 ;
      RECT  7.165 2.92 7.395 3.245 ;
      RECT  6.045 3.245 7.395 3.475 ;
      RECT  6.045 3.475 6.275 3.805 ;
      RECT  0.18 3.805 6.275 4.035 ;
      RECT  7.67 4.985 12.49 5.215 ;
  END
END MDN_AN3B_3
#-----------------------------------------------------------------------
#      Cell        : MDN_AN3B_4
#      Description : 3-Input AND (A inverted input)
#      Equation    : X=!A&B1&B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN3B_4
  CLASS CORE ;
  FOREIGN MDN_AN3B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.93 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.93 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  7.725 4.93 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.695 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.695 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  12.205 0.14 12.435 0.695 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.63 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.685 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.13 1.005 17.74 1.235 ;
      RECT  13.325 1.235 13.555 3.245 ;
      RECT  9.965 3.245 13.555 3.475 ;
      RECT  9.965 3.475 10.195 3.805 ;
      RECT  9.13 3.805 10.195 4.035 ;
    END
    ANTENNADIFFAREA 8.18 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 8.78 1.235 ;
      RECT  5.43 1.565 9.635 1.795 ;
      RECT  9.405 1.795 9.635 2.405 ;
      RECT  9.405 2.405 12.945 2.635 ;
      RECT  9.405 2.635 9.635 3.245 ;
      RECT  8.285 3.245 9.635 3.475 ;
      RECT  8.285 3.475 8.515 4.365 ;
      RECT  0.18 4.365 8.515 4.595 ;
      RECT  11.085 4.365 17.74 4.595 ;
      RECT  11.085 4.595 11.315 4.925 ;
      RECT  9.895 4.925 11.315 5.155 ;
  END
END MDN_AN3B_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AN4_1
#      Description : 4-Input AND
#      Equation    : X=A1&A2&A3&A4
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN4_1
  CLASS CORE ;
  FOREIGN MDN_AN4_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  1.005 5.46 3.475 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 3.245 ;
      RECT  4.66 3.245 5.155 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  4.365 0.37 5.21 0.6 ;
      RECT  4.365 0.6 4.595 1.005 ;
      RECT  3.245 1.005 4.595 1.235 ;
      RECT  3.245 1.235 3.475 4.365 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  1.72 1.005 2.76 1.235 ;
  END
END MDN_AN4_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AN4_2
#      Description : 4-Input AND
#      Equation    : X=A1&A2&A3&A4
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN4_2
  CLASS CORE ;
  FOREIGN MDN_AN4_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  3.245 5.46 5.715 5.74 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  0.56 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 6.54 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  4.66 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  3.245 1.005 4.3 1.235 ;
      RECT  3.245 1.235 3.475 4.365 ;
      RECT  0.18 4.365 6.22 4.595 ;
      RECT  4.98 4.595 5.21 5.0 ;
      RECT  5.99 4.595 6.22 5.0 ;
      RECT  4.87 5.0 5.21 5.23 ;
      RECT  5.99 5.0 6.33 5.23 ;
  END
END MDN_AN4_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AN4_4
#      Description : 4-Input AND
#      Equation    : X=A1&A2&A3&A4
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN4_4
  CLASS CORE ;
  FOREIGN MDN_AN4_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.93 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  1.005 5.46 3.475 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  0.0 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 8.78 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  4.66 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 8.57 0.6 ;
      RECT  8.23 0.6 8.46 1.005 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  7.22 0.6 7.45 1.005 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  3.245 1.005 6.22 1.235 ;
      RECT  7.22 1.005 8.46 1.235 ;
      RECT  3.245 1.235 3.475 4.365 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  1.72 1.005 2.76 1.235 ;
  END
END MDN_AN4_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AN4B_1
#      Description : 4-Input AND (A inverted input)
#      Equation    : X=!A&B1&B2&B3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN4B_1
  CLASS CORE ;
  FOREIGN MDN_AN4B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 4.365 6.54 4.595 ;
      RECT  6.045 4.595 6.275 5.46 ;
      RECT  6.045 5.46 6.89 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  1.005 5.46 1.68 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  4.31 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  1.005 -0.14 1.68 0.14 ;
      RECT  1.005 0.14 1.235 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.005 6.54 1.235 ;
      RECT  4.925 1.235 5.155 4.365 ;
      RECT  4.66 4.365 5.155 4.595 ;
    END
    ANTENNADIFFAREA 2.126 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.805 0.37 5.21 0.6 ;
      RECT  3.805 0.6 4.035 1.565 ;
      RECT  3.805 1.565 4.595 1.795 ;
      RECT  4.365 1.795 4.595 3.805 ;
      RECT  3.805 3.805 4.595 4.035 ;
      RECT  3.805 4.035 4.035 4.365 ;
      RECT  1.72 4.365 4.035 4.595 ;
      RECT  1.72 1.005 2.76 1.235 ;
  END
END MDN_AN4B_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AN4B_2
#      Description : 4-Input AND (A inverted input)
#      Equation    : X=!A&B1&B2&B3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN4B_2
  CLASS CORE ;
  FOREIGN MDN_AN4B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.905 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  3.245 5.46 4.65 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  1.005 5.46 1.68 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  1.005 -0.14 2.41 0.14 ;
      RECT  1.005 0.14 1.235 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.005 8.78 1.235 ;
      RECT  4.91 1.235 5.14 3.245 ;
      RECT  4.91 3.245 5.77 3.475 ;
    END
    ANTENNADIFFAREA 3.928 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  3.96 1.565 4.595 1.795 ;
      RECT  4.365 1.795 4.595 3.805 ;
      RECT  3.805 3.805 4.595 4.035 ;
      RECT  3.805 4.035 4.035 4.365 ;
      RECT  1.72 4.365 4.035 4.595 ;
      RECT  3.805 4.595 4.035 4.995 ;
      RECT  3.805 4.995 6.14 5.0 ;
      RECT  3.805 5.0 6.33 5.23 ;
      RECT  4.66 4.365 8.78 4.595 ;
  END
END MDN_AN4B_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AN4B_3
#      Description : 4-Input AND (A inverted input)
#      Equation    : X=!A&B1&B2&B3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN4B_3
  CLASS CORE ;
  FOREIGN MDN_AN4B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.115 10.715 2.125 ;
      RECT  8.26 2.125 10.78 2.345 ;
      RECT  8.26 2.345 8.54 2.915 ;
      RECT  9.38 2.345 9.66 2.915 ;
      RECT  10.5 2.345 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.74 0.37 4.08 0.6 ;
      RECT  3.78 0.6 4.06 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  8.44 4.365 11.02 4.595 ;
      RECT  10.525 4.595 10.755 5.46 ;
      RECT  10.08 5.46 11.37 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.595 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.595 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 1.005 11.02 1.235 ;
      RECT  7.725 1.235 7.955 1.565 ;
      RECT  4.66 1.565 7.955 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  4.66 3.245 7.955 3.475 ;
    END
    ANTENNADIFFAREA 6.378 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  3.805 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 2.405 ;
      RECT  3.805 2.405 7.39 2.635 ;
      RECT  3.805 2.635 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
      RECT  3.805 3.475 4.035 3.805 ;
      RECT  1.72 3.805 4.035 4.035 ;
      RECT  5.43 4.925 10.25 5.155 ;
  END
END MDN_AN4B_3
#-----------------------------------------------------------------------
#      Cell        : MDN_AN4B_4
#      Description : 4-Input AND (A inverted input)
#      Equation    : X=!A&B1&B2&B3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AN4B_4
  CLASS CORE ;
  FOREIGN MDN_AN4B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.39 2.115 12.955 2.125 ;
      RECT  9.38 2.125 13.02 2.345 ;
      RECT  9.38 2.345 9.66 2.915 ;
      RECT  10.5 2.345 10.78 2.915 ;
      RECT  11.62 2.345 11.9 2.915 ;
      RECT  12.74 2.345 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.75 0.37 4.09 0.6 ;
      RECT  3.78 0.6 4.06 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.93 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.93 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.905 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.695 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.845 1.005 13.26 1.235 ;
      RECT  8.845 1.235 9.075 1.565 ;
      RECT  4.66 1.565 9.075 1.795 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  4.66 3.245 9.075 3.475 ;
    END
    ANTENNADIFFAREA 8.504 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  3.805 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 2.405 ;
      RECT  3.805 2.405 8.48 2.635 ;
      RECT  3.805 2.635 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
      RECT  3.805 3.475 4.035 3.805 ;
      RECT  1.72 3.805 4.035 4.035 ;
      RECT  8.845 4.365 13.26 4.595 ;
      RECT  8.845 4.595 9.075 4.925 ;
      RECT  5.43 4.925 9.075 5.155 ;
  END
END MDN_AN4B_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AO2111_1
#      Description : One 2-input AND into 4-input OR
#      Equation    : X=(A1&A2)|B1|B2|B3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO2111_1
  CLASS CORE ;
  FOREIGN MDN_AO2111_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 7.42 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 8.54 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 4.365 4.06 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.93 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.925 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.925 1.235 5.46 ;
      RECT  1.005 5.46 2.41 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  8.285 -0.14 8.96 0.14 ;
      RECT  8.285 0.14 8.515 1.005 ;
      RECT  8.285 1.005 8.78 1.235 ;
      RECT  3.245 -0.14 5.155 0.14 ;
      RECT  3.245 0.14 3.475 0.585 ;
      RECT  4.925 0.14 5.155 1.005 ;
      RECT  4.66 1.005 5.155 1.235 ;
      RECT  1.005 -0.14 1.68 0.14 ;
      RECT  1.005 0.14 1.235 0.585 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 1.005 6.54 1.235 ;
      RECT  5.485 1.235 5.715 3.245 ;
      RECT  4.62 3.245 5.715 3.475 ;
      RECT  5.485 3.475 5.715 4.365 ;
      RECT  5.485 4.365 6.54 4.595 ;
    END
    ANTENNADIFFAREA 2.41 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.67 1.005 4.3 1.235 ;
      RECT  3.805 1.235 4.035 2.38 ;
      RECT  3.805 2.38 5.065 2.61 ;
      RECT  3.805 2.61 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
      RECT  6.045 1.565 7.24 1.795 ;
      RECT  6.045 1.795 6.275 3.805 ;
      RECT  6.045 3.805 7.395 4.035 ;
      RECT  7.165 4.035 7.395 4.365 ;
      RECT  7.165 4.365 8.78 4.595 ;
      RECT  1.67 4.365 2.76 4.595 ;
  END
END MDN_AO2111_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AO2111_2
#      Description : One 2-input AND into 4-input OR
#      Equation    : X=(A1&A2)|B1|B2|B3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO2111_2
  CLASS CORE ;
  FOREIGN MDN_AO2111_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 4.365 4.06 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.925 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.925 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.925 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.925 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.525 -0.14 11.37 0.14 ;
      RECT  10.525 0.14 10.755 1.005 ;
      RECT  10.525 1.005 11.02 1.235 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 1.005 8.78 1.235 ;
      RECT  7.725 1.235 7.955 1.565 ;
      RECT  6.605 1.565 7.955 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  4.62 3.245 7.955 3.475 ;
      RECT  7.725 3.475 7.955 3.805 ;
      RECT  7.725 3.805 8.885 4.035 ;
    END
    ANTENNADIFFAREA 4.82 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  7.165 0.445 8.01 0.675 ;
      RECT  7.165 0.675 7.395 1.005 ;
      RECT  4.62 1.005 7.395 1.235 ;
      RECT  1.67 1.005 4.3 1.235 ;
      RECT  3.805 1.235 4.035 2.405 ;
      RECT  3.805 2.405 6.33 2.635 ;
      RECT  3.805 2.635 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
      RECT  8.285 1.565 9.48 1.795 ;
      RECT  8.285 1.795 8.515 2.405 ;
      RECT  7.11 2.405 8.515 2.635 ;
      RECT  8.285 2.635 8.515 3.245 ;
      RECT  8.285 3.245 9.635 3.475 ;
      RECT  9.405 3.475 9.635 3.805 ;
      RECT  9.405 3.805 11.02 4.035 ;
      RECT  1.67 4.365 2.76 4.595 ;
  END
END MDN_AO2111_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AO2111_4
#      Description : One 2-input AND into 4-input OR
#      Equation    : X=(A1&A2)|B1|B2|B3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO2111_4
  CLASS CORE ;
  FOREIGN MDN_AO2111_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 14.14 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.98 2.125 15.26 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 4.365 4.06 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.925 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.925 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.965 4.925 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.925 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.925 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.925 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  15.005 -0.14 15.85 0.14 ;
      RECT  15.005 0.14 15.235 1.005 ;
      RECT  15.005 1.005 15.5 1.235 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 1.005 13.26 1.235 ;
      RECT  12.205 1.235 12.435 1.565 ;
      RECT  8.845 1.565 12.435 1.795 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  4.62 3.245 12.435 3.475 ;
      RECT  12.205 3.475 12.435 3.805 ;
      RECT  12.205 3.805 13.26 4.035 ;
    END
    ANTENNADIFFAREA 9.64 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.845 0.445 12.49 0.675 ;
      RECT  8.845 0.675 9.075 1.005 ;
      RECT  8.285 1.005 9.075 1.235 ;
      RECT  8.285 1.235 8.515 1.565 ;
      RECT  4.62 1.565 8.515 1.795 ;
      RECT  1.67 1.005 4.3 1.235 ;
      RECT  3.805 1.235 4.035 2.405 ;
      RECT  3.805 2.405 8.58 2.635 ;
      RECT  3.805 2.635 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
      RECT  12.765 1.565 13.96 1.795 ;
      RECT  12.765 1.795 12.995 2.405 ;
      RECT  9.35 2.405 12.995 2.635 ;
      RECT  12.765 2.635 12.995 3.245 ;
      RECT  12.765 3.245 14.115 3.475 ;
      RECT  13.885 3.475 14.115 3.805 ;
      RECT  13.885 3.805 15.5 4.035 ;
      RECT  1.67 4.365 2.76 4.595 ;
  END
END MDN_AO2111_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AO211_1
#      Description : One 2-input AND into 3-input OR
#      Equation    : X=(A1&A2)|B1|B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO211_1
  CLASS CORE ;
  FOREIGN MDN_AO211_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 4.365 4.06 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  0.0 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 3.245 ;
      RECT  4.66 3.245 5.155 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  4.365 0.37 5.21 0.6 ;
      RECT  4.365 0.6 4.595 1.005 ;
      RECT  1.72 1.005 4.595 1.235 ;
      RECT  3.805 1.235 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
      RECT  0.18 4.365 2.76 4.595 ;
  END
END MDN_AO211_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AO211_2
#      Description : One 2-input AND into 3-input OR
#      Equation    : X=(A1&A2)|B1|B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO211_2
  CLASS CORE ;
  FOREIGN MDN_AO211_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 4.365 4.06 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 6.89 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  0.0 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 6.54 1.795 ;
      RECT  4.925 1.795 5.155 3.245 ;
      RECT  4.66 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  1.72 1.005 6.22 1.235 ;
      RECT  3.805 1.235 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
      RECT  0.18 4.365 2.76 4.595 ;
  END
END MDN_AO211_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AO211_4
#      Description : One 2-input AND into 3-input OR
#      Equation    : X=(A1&A2)|B1|B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO211_4
  CLASS CORE ;
  FOREIGN MDN_AO211_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 4.365 4.06 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.93 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  0.0 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 8.78 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  4.66 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 8.57 0.6 ;
      RECT  8.23 0.6 8.46 1.005 ;
      RECT  5.97 0.37 7.45 0.6 ;
      RECT  7.22 0.6 7.45 1.005 ;
      RECT  7.22 1.005 8.46 1.235 ;
      RECT  1.72 1.005 4.035 1.235 ;
      RECT  3.805 1.235 4.035 1.565 ;
      RECT  3.805 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 2.405 ;
      RECT  3.805 2.405 6.33 2.635 ;
      RECT  3.805 2.635 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
      RECT  0.18 4.365 2.76 4.595 ;
  END
END MDN_AO211_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AO21_1
#      Description : One 2-input AND into 2-input OR
#      Equation    : X=(A1&A2)|B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO21_1
  CLASS CORE ;
  FOREIGN MDN_AO21_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.445 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.745 0.37 4.09 0.6 ;
      RECT  3.745 0.6 3.975 1.005 ;
      RECT  1.005 0.445 2.915 0.675 ;
      RECT  2.685 0.675 2.915 1.005 ;
      RECT  1.005 0.675 1.235 3.805 ;
      RECT  2.685 1.005 3.975 1.235 ;
      RECT  0.16 3.805 1.235 4.035 ;
      RECT  1.675 1.005 2.355 1.235 ;
      RECT  2.125 1.235 2.355 1.565 ;
      RECT  2.125 1.565 2.76 1.795 ;
      RECT  2.475 4.34 2.705 4.925 ;
      RECT  0.905 4.925 2.705 5.155 ;
  END
END MDN_AO21_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AO21_2
#      Description : One 2-input AND into 2-input OR
#      Equation    : X=(A1&A2)|B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO21_2
  CLASS CORE ;
  FOREIGN MDN_AO21_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.445 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  0.0 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  3.96 3.245 5.0 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  3.75 0.6 3.98 1.005 ;
      RECT  1.005 0.445 2.9 0.675 ;
      RECT  2.67 0.675 2.9 1.005 ;
      RECT  1.005 0.675 1.235 3.805 ;
      RECT  2.67 1.005 3.98 1.235 ;
      RECT  0.18 3.805 1.235 4.035 ;
      RECT  1.675 1.005 2.355 1.235 ;
      RECT  2.125 1.235 2.355 1.565 ;
      RECT  2.125 1.565 2.76 1.795 ;
      RECT  2.475 4.34 2.705 4.925 ;
      RECT  0.95 4.925 2.705 5.155 ;
  END
END MDN_AO21_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AO21_3
#      Description : One 2-input AND into 2-input OR
#      Equation    : X=(A1&A2)|B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO21_3
  CLASS CORE ;
  FOREIGN MDN_AO21_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.445 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  0.0 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.96 1.565 6.54 1.795 ;
      RECT  4.92 1.795 5.15 3.245 ;
      RECT  3.765 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 4.536 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  3.75 0.6 3.98 1.005 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  1.005 0.445 2.915 0.675 ;
      RECT  2.685 0.675 2.915 1.005 ;
      RECT  1.005 0.675 1.235 3.805 ;
      RECT  2.685 1.005 3.98 1.235 ;
      RECT  4.98 1.005 6.22 1.235 ;
      RECT  0.16 3.805 1.235 4.035 ;
      RECT  1.675 1.005 2.355 1.235 ;
      RECT  2.125 1.235 2.355 1.565 ;
      RECT  2.125 1.565 2.76 1.795 ;
      RECT  2.475 4.34 2.705 4.925 ;
      RECT  0.905 4.925 2.705 5.155 ;
  END
END MDN_AO21_3
#-----------------------------------------------------------------------
#      Cell        : MDN_AO21_4
#      Description : One 2-input AND into 2-input OR
#      Equation    : X=(A1&A2)|B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO21_4
  CLASS CORE ;
  FOREIGN MDN_AO21_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  0.445 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.765 1.565 7.38 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  3.765 3.245 7.38 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  3.75 0.6 3.98 1.005 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  1.005 0.445 2.9 0.675 ;
      RECT  2.67 0.675 2.9 1.005 ;
      RECT  1.005 0.675 1.235 3.805 ;
      RECT  2.67 1.005 3.98 1.235 ;
      RECT  4.98 1.005 6.22 1.235 ;
      RECT  0.16 3.805 1.235 4.035 ;
      RECT  1.675 1.005 2.355 1.235 ;
      RECT  2.125 1.235 2.355 1.565 ;
      RECT  2.125 1.565 2.76 1.795 ;
      RECT  2.475 4.34 2.705 4.925 ;
      RECT  0.95 4.925 2.705 5.155 ;
  END
END MDN_AO21_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AO21_6
#      Description : One 2-input AND into 2-input OR
#      Equation    : X=(A1&A2)|B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO21_6
  CLASS CORE ;
  FOREIGN MDN_AO21_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.685 ;
      RECT  2.66 2.685 4.06 2.915 ;
      RECT  3.78 2.125 4.06 2.685 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.905 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.905 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 4.905 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.695 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.005 7.395 1.235 ;
      RECT  7.165 1.235 7.395 1.565 ;
      RECT  7.165 1.565 13.26 1.795 ;
      RECT  11.085 1.795 11.315 3.245 ;
      RECT  7.165 3.245 13.26 3.475 ;
      RECT  7.165 3.475 7.395 4.365 ;
      RECT  6.9 4.365 7.395 4.595 ;
    END
    ANTENNADIFFAREA 9.072 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 11.93 0.6 ;
      RECT  3.19 0.445 4.945 0.675 ;
      RECT  4.715 0.675 4.945 1.005 ;
      RECT  4.715 1.005 6.275 1.235 ;
      RECT  6.045 1.235 6.275 1.565 ;
      RECT  6.045 1.565 6.835 1.795 ;
      RECT  6.605 1.795 6.835 2.125 ;
      RECT  6.605 2.125 10.755 2.355 ;
      RECT  7.165 2.355 7.395 2.69 ;
      RECT  8.285 2.355 8.515 2.69 ;
      RECT  9.405 2.355 9.635 2.69 ;
      RECT  10.525 2.355 10.755 2.69 ;
      RECT  6.605 2.355 6.835 3.805 ;
      RECT  6.045 3.805 6.835 4.035 ;
      RECT  6.045 4.035 6.275 4.365 ;
      RECT  4.64 4.365 6.275 4.595 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  11.645 2.125 12.995 2.355 ;
      RECT  11.645 2.355 11.875 2.69 ;
      RECT  12.765 2.355 12.995 2.69 ;
      RECT  0.175 4.365 4.3 4.595 ;
      RECT  4.07 4.595 4.3 4.925 ;
      RECT  4.07 4.925 5.77 5.155 ;
  END
END MDN_AO21_6
#-----------------------------------------------------------------------
#      Cell        : MDN_AO21B_1
#      Description : One 2-input NAND into 2-input NAND
#      Equation    : X=(A1&A2)|!B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO21B_1
  CLASS CORE ;
  FOREIGN MDN_AO21B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 4.48 5.74 ;
      RECT  1.72 4.365 2.76 4.595 ;
      RECT  2.125 4.595 2.355 5.46 ;
      RECT  1.68 5.46 2.8 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  0.0 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 -0.14 4.48 0.14 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  2.685 1.235 2.915 3.245 ;
      RECT  2.685 3.245 3.53 3.475 ;
    END
    ANTENNADIFFAREA 2.086 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.83 0.37 2.99 0.6 ;
      RECT  1.83 0.6 2.06 1.005 ;
      RECT  1.005 1.005 2.06 1.235 ;
      RECT  1.005 1.235 1.235 3.475 ;
  END
END MDN_AO21B_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AO21B_2
#      Description : One 2-input NAND into 2-input NAND
#      Equation    : X=(A1&A2)|!B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO21B_2
  CLASS CORE ;
  FOREIGN MDN_AO21B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  1.005 5.46 3.475 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 4.595 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  2.42 3.245 4.595 3.475 ;
      RECT  4.365 3.475 4.595 3.805 ;
      RECT  4.365 3.805 6.54 4.035 ;
    END
    ANTENNADIFFAREA 4.82 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.445 4.595 0.675 ;
      RECT  4.365 0.675 4.595 1.005 ;
      RECT  4.365 1.005 6.54 1.235 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.395 ;
      RECT  1.565 2.395 4.09 2.625 ;
      RECT  1.565 2.625 1.795 3.805 ;
      RECT  0.18 3.805 2.06 4.035 ;
  END
END MDN_AO21B_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AO21B_3
#      Description : One 2-input NAND into 2-input NAND
#      Equation    : X=(A1&A2)|!B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO21B_3
  CLASS CORE ;
  FOREIGN MDN_AO21B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 8.54 2.355 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 5.715 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  0.56 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.84 -0.14 9.13 0.14 ;
      RECT  8.285 0.14 8.515 1.005 ;
      RECT  6.2 1.005 8.78 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 5.0 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  2.42 3.245 4.595 3.475 ;
      RECT  4.365 3.475 4.595 3.805 ;
      RECT  4.365 3.805 8.78 4.035 ;
    END
    ANTENNADIFFAREA 7.23 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.445 8.01 0.675 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.41 ;
      RECT  1.565 2.41 4.09 2.64 ;
      RECT  1.565 2.64 1.795 3.805 ;
      RECT  0.18 3.805 2.06 4.035 ;
      RECT  3.75 5.0 5.21 5.23 ;
  END
END MDN_AO21B_3
#-----------------------------------------------------------------------
#      Cell        : MDN_AO21B_4
#      Description : One 2-input NAND into 2-input NAND
#      Equation    : X=(A1&A2)|!B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO21B_4
  CLASS CORE ;
  FOREIGN MDN_AO21B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.54 0.6 1.82 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 10.78 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 5.715 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 6.54 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  2.42 3.245 4.595 3.475 ;
      RECT  4.365 3.475 4.595 3.805 ;
      RECT  4.365 3.805 11.02 4.035 ;
    END
    ANTENNADIFFAREA 9.64 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.445 6.835 0.675 ;
      RECT  6.605 0.675 6.835 1.005 ;
      RECT  6.605 1.005 11.02 1.235 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.4 ;
      RECT  1.565 2.4 4.09 2.63 ;
      RECT  1.565 2.63 1.795 3.805 ;
      RECT  0.18 3.805 2.06 4.035 ;
      RECT  4.87 2.4 6.33 2.63 ;
      RECT  3.75 5.0 5.21 5.23 ;
  END
END MDN_AO21B_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AO221_1
#      Description : Two 2-input ANDs into 3 input OR
#      Equation    : X=(A1&A2)|(B1&B2)|C
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO221_1
  CLASS CORE ;
  FOREIGN MDN_AO221_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.36 5.46 4.035 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.725 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.95 0.37 6.33 0.6 ;
      RECT  5.95 0.6 6.18 1.005 ;
      RECT  3.245 0.445 5.155 0.675 ;
      RECT  4.925 0.675 5.155 1.005 ;
      RECT  3.245 0.675 3.475 1.565 ;
      RECT  4.925 1.005 6.18 1.235 ;
      RECT  1.72 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 3.245 ;
      RECT  2.685 3.245 3.475 3.475 ;
      RECT  2.685 3.475 2.915 3.805 ;
      RECT  1.72 3.805 2.915 4.035 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.005 4.595 1.235 ;
      RECT  4.365 1.235 4.595 1.565 ;
      RECT  4.365 1.565 5.0 1.795 ;
      RECT  3.245 3.805 5.0 4.035 ;
      RECT  3.245 4.035 3.475 4.925 ;
      RECT  0.235 4.31 0.465 4.925 ;
      RECT  0.235 4.925 3.475 5.155 ;
      RECT  0.95 4.365 2.76 4.595 ;
  END
END MDN_AO221_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AO221_2
#      Description : Two 2-input ANDs into 3 input OR
#      Equation    : X=(A1&A2)|(B1&B2)|C
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO221_2
  CLASS CORE ;
  FOREIGN MDN_AO221_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 9.13 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.36 5.46 4.035 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.735 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 7.395 1.795 ;
      RECT  7.165 1.795 7.395 3.245 ;
      RECT  6.2 3.245 7.395 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.245 0.445 5.155 0.675 ;
      RECT  4.925 0.675 5.155 1.005 ;
      RECT  3.245 0.675 3.475 1.565 ;
      RECT  4.925 1.005 6.22 1.235 ;
      RECT  1.72 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 3.245 ;
      RECT  2.685 3.245 3.475 3.475 ;
      RECT  2.685 3.475 2.915 3.805 ;
      RECT  1.72 3.805 2.915 4.035 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.005 4.595 1.235 ;
      RECT  4.365 1.235 4.595 1.565 ;
      RECT  4.365 1.565 5.0 1.795 ;
      RECT  3.245 3.805 5.0 4.035 ;
      RECT  3.245 4.035 3.475 4.925 ;
      RECT  0.235 4.31 0.465 4.925 ;
      RECT  0.235 4.925 3.475 5.155 ;
      RECT  0.95 4.365 2.76 4.595 ;
  END
END MDN_AO221_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AO221_4
#      Description : Two 2-input ANDs into 3 input OR
#      Equation    : X=(A1&A2)|(B1&B2)|C
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO221_4
  CLASS CORE ;
  FOREIGN MDN_AO221_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.36 5.46 4.035 5.74 ;
      RECT  -0.17 5.46 0.56 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 9.485 1.795 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  6.2 3.245 9.48 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 9.69 0.6 ;
      RECT  3.245 0.445 5.155 0.675 ;
      RECT  4.925 0.675 5.155 1.005 ;
      RECT  3.245 0.675 3.475 1.565 ;
      RECT  4.925 1.005 5.715 1.235 ;
      RECT  5.485 1.235 5.715 2.125 ;
      RECT  1.72 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 3.245 ;
      RECT  5.485 2.125 8.515 2.355 ;
      RECT  6.045 2.355 6.275 2.69 ;
      RECT  7.165 2.355 7.395 2.69 ;
      RECT  8.285 2.355 8.515 2.69 ;
      RECT  2.685 3.245 3.475 3.475 ;
      RECT  2.685 3.475 2.915 3.805 ;
      RECT  1.72 3.805 2.915 4.035 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.005 4.595 1.235 ;
      RECT  4.365 1.235 4.595 1.565 ;
      RECT  4.365 1.565 5.0 1.795 ;
      RECT  3.245 3.805 5.0 4.035 ;
      RECT  3.245 4.035 3.475 4.925 ;
      RECT  0.235 4.34 0.465 4.925 ;
      RECT  0.235 4.925 3.475 5.155 ;
      RECT  0.95 4.365 2.76 4.595 ;
  END
END MDN_AO221_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AO22_1
#      Description : Two 2-input ANDs into 2-input OR
#      Equation    : X=(A1&A2)|(B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO22_1
  CLASS CORE ;
  FOREIGN MDN_AO22_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  1.005 5.46 2.41 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  4.31 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 1.005 ;
      RECT  3.96 1.005 5.715 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 3.245 ;
      RECT  4.66 3.245 5.155 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.245 0.37 5.21 0.6 ;
      RECT  3.245 0.6 3.475 1.005 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 3.5 ;
      RECT  0.18 4.365 4.3 4.595 ;
  END
END MDN_AO22_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AO22_2
#      Description : Two 2-input ANDs into 2-input OR
#      Equation    : X=(A1&A2)|(B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO22_2
  CLASS CORE ;
  FOREIGN MDN_AO22_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 6.54 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  4.66 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 4.365 ;
      RECT  2.42 4.365 6.22 4.595 ;
      RECT  4.98 4.595 5.21 5.0 ;
      RECT  5.99 4.595 6.22 5.0 ;
      RECT  4.87 5.0 5.21 5.23 ;
      RECT  5.99 5.0 6.33 5.23 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  1.83 4.595 2.06 4.925 ;
      RECT  1.83 4.925 3.53 5.155 ;
  END
END MDN_AO22_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AO22_3
#      Description : Two 2-input ANDs into 2-input OR
#      Equation    : X=(A1&A2)|(B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO22_3
  CLASS CORE ;
  FOREIGN MDN_AO22_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  3.36 -0.14 4.035 0.14 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.005 5.715 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  5.485 1.565 7.24 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  4.66 3.245 7.24 3.475 ;
    END
    ANTENNADIFFAREA 4.536 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.98 0.37 7.45 0.6 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  3.245 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 2.685 ;
      RECT  4.925 2.685 6.275 2.915 ;
      RECT  6.045 2.35 6.275 2.685 ;
      RECT  2.42 4.365 4.3 4.595 ;
      RECT  4.07 4.595 4.3 5.0 ;
      RECT  4.07 5.0 5.19 5.23 ;
      RECT  0.95 4.925 3.53 5.155 ;
  END
END MDN_AO22_3
#-----------------------------------------------------------------------
#      Cell        : MDN_AO22_4
#      Description : Two 2-input ANDs into 2-input OR
#      Equation    : X=(A1&A2)|(B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO22_4
  CLASS CORE ;
  FOREIGN MDN_AO22_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  1.005 5.46 2.41 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  3.805 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.005 5.715 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  5.485 1.565 8.78 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  4.66 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 8.57 0.6 ;
      RECT  8.23 0.6 8.46 1.005 ;
      RECT  7.095 0.37 7.45 0.6 ;
      RECT  7.22 0.6 7.45 1.005 ;
      RECT  7.22 1.005 8.46 1.235 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  3.245 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 2.125 ;
      RECT  3.245 1.795 3.475 3.5 ;
      RECT  4.925 2.125 7.395 2.355 ;
      RECT  4.925 2.355 5.155 2.69 ;
      RECT  6.045 2.355 6.275 2.69 ;
      RECT  7.165 2.355 7.395 2.69 ;
      RECT  0.18 4.365 4.3 4.595 ;
  END
END MDN_AO22_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AO22_6
#      Description : Two 2-input ANDs into 2-input OR
#      Equation    : X=(A1&A2)|(B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO22_6
  CLASS CORE ;
  FOREIGN MDN_AO22_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.14 1.565 15.5 1.795 ;
      RECT  13.325 1.795 13.555 3.245 ;
      RECT  9.14 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 9.072 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  14.95 0.37 15.29 0.6 ;
      RECT  14.95 0.6 15.18 1.005 ;
      RECT  12.71 0.37 14.17 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  13.94 0.6 14.17 1.005 ;
      RECT  10.47 0.37 11.93 0.6 ;
      RECT  10.47 0.6 10.7 1.005 ;
      RECT  11.7 0.6 11.93 1.005 ;
      RECT  9.35 0.37 9.69 0.6 ;
      RECT  9.46 0.6 9.69 1.005 ;
      RECT  7.15 1.005 10.7 1.235 ;
      RECT  11.7 1.005 12.94 1.235 ;
      RECT  13.94 1.005 15.18 1.235 ;
      RECT  7.15 1.235 7.38 1.565 ;
      RECT  2.42 1.005 4.035 1.235 ;
      RECT  3.805 1.235 4.035 1.565 ;
      RECT  3.805 1.565 7.38 1.795 ;
      RECT  6.605 1.795 6.835 4.365 ;
      RECT  4.66 4.365 8.78 4.595 ;
      RECT  1.83 0.445 3.53 0.675 ;
      RECT  1.83 0.675 2.06 1.005 ;
      RECT  0.18 1.005 2.06 1.235 ;
      RECT  6.605 0.445 8.01 0.675 ;
      RECT  6.605 0.675 6.835 1.005 ;
      RECT  4.66 1.005 6.835 1.235 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.07 4.595 4.3 4.925 ;
      RECT  4.07 4.925 8.01 5.155 ;
  END
END MDN_AO22_6
#-----------------------------------------------------------------------
#      Cell        : MDN_AO2BB2_1
#      Description : One 2-input AND with inverted inputs + 2-input AND into 2-input OR
#      Equation    : X=(!A1&!A2)|(B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO2BB2_1
  CLASS CORE ;
  FOREIGN MDN_AO2BB2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  2.42 4.365 2.915 4.595 ;
      RECT  2.685 4.595 2.915 5.46 ;
      RECT  2.24 5.46 2.915 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 1.565 ;
      RECT  3.96 1.565 5.715 1.795 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 3.53 ;
    END
    ANTENNADIFFAREA 2.086 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.445 4.595 0.675 ;
      RECT  4.365 0.675 4.595 1.005 ;
      RECT  4.365 1.005 5.0 1.235 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.805 ;
      RECT  1.83 3.805 2.915 4.035 ;
      RECT  1.83 4.035 2.06 4.365 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  3.96 4.365 5.0 4.595 ;
  END
END MDN_AO2BB2_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AO2BB2_2
#      Description : One 2-input AND with inverted inputs + 2-input AND into 2-input OR
#      Equation    : X=(!A1&!A2)|(B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO2BB2_2
  CLASS CORE ;
  FOREIGN MDN_AO2BB2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 1.51 3.475 4.365 ;
      RECT  2.42 4.365 6.54 4.595 ;
    END
    ANTENNADIFFAREA 4.686 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  2.63 0.37 4.09 0.6 ;
      RECT  2.42 1.005 8.78 1.235 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.805 ;
      RECT  1.565 3.805 2.915 4.035 ;
      RECT  1.565 4.035 1.795 4.365 ;
      RECT  0.18 4.365 1.795 4.595 ;
      RECT  6.9 4.365 8.78 4.595 ;
      RECT  6.9 4.595 7.13 4.925 ;
      RECT  5.43 4.925 7.13 5.155 ;
  END
END MDN_AO2BB2_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AO2BB2_4
#      Description : One 2-input AND with inverted inputs + 2-input AND into 2-input OR
#      Equation    : X=(!A1&!A2)|(B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO2BB2_4
  CLASS CORE ;
  FOREIGN MDN_AO2BB2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 10.78 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 2.125 15.26 2.355 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.87 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.905 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.19 1.565 5.77 1.795 ;
      RECT  4.365 1.795 4.595 4.365 ;
      RECT  2.42 4.365 11.02 4.595 ;
    END
    ANTENNADIFFAREA 9.372 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 6.33 0.6 ;
      RECT  2.42 1.005 15.5 1.235 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 2.405 ;
      RECT  2.685 2.405 4.09 2.635 ;
      RECT  2.685 2.635 2.915 3.805 ;
      RECT  1.565 3.805 2.915 4.035 ;
      RECT  1.565 4.035 1.795 4.365 ;
      RECT  0.14 4.365 1.795 4.595 ;
      RECT  11.34 4.365 15.5 4.595 ;
      RECT  11.34 4.595 11.57 4.925 ;
      RECT  7.67 4.925 11.57 5.155 ;
  END
END MDN_AO2BB2_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AO311_1
#      Description : One 3-input AND into 3-input OR
#      Equation    : X=(A1&A2&A3)|B1|B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO311_1
  CLASS CORE ;
  FOREIGN MDN_AO311_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 6.89 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.95 0.37 6.33 0.6 ;
      RECT  5.95 0.6 6.18 1.005 ;
      RECT  5.49 1.005 6.18 1.235 ;
      RECT  5.49 1.235 5.72 1.565 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 1.565 ;
      RECT  1.005 1.565 5.72 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  3.96 3.245 4.595 3.475 ;
      RECT  1.72 1.005 5.0 1.235 ;
      RECT  4.365 4.365 5.0 4.595 ;
      RECT  4.365 4.595 4.595 4.925 ;
      RECT  0.18 4.365 2.915 4.595 ;
      RECT  2.685 4.595 2.915 4.925 ;
      RECT  2.685 4.925 4.595 5.155 ;
  END
END MDN_AO311_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AO311_2
#      Description : One 3-input AND into 3-input OR
#      Equation    : X=(A1&A2&A3)|B1|B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO311_2
  CLASS CORE ;
  FOREIGN MDN_AO311_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.905 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.905 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  6.2 3.245 7.24 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  5.485 1.005 6.22 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 1.565 ;
      RECT  1.005 1.565 5.715 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  3.96 3.245 4.595 3.475 ;
      RECT  1.72 1.005 5.0 1.235 ;
      RECT  4.365 4.365 5.0 4.595 ;
      RECT  4.365 4.595 4.595 4.925 ;
      RECT  0.18 4.365 2.915 4.595 ;
      RECT  2.685 4.595 2.915 4.925 ;
      RECT  2.685 4.925 4.595 5.155 ;
  END
END MDN_AO311_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AO311_4
#      Description : One 3-input AND into 3-input OR
#      Equation    : X=(A1&A2&A3)|B1|B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO311_4
  CLASS CORE ;
  FOREIGN MDN_AO311_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 11.37 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 9.48 1.795 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  6.2 3.245 9.48 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.22 0.37 9.69 0.6 ;
      RECT  0.14 1.005 5.0 1.235 ;
      RECT  1.67 1.565 5.715 1.795 ;
      RECT  5.485 1.795 5.715 2.125 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  5.485 2.125 8.515 2.355 ;
      RECT  6.045 2.355 6.275 2.69 ;
      RECT  7.165 2.355 7.395 2.69 ;
      RECT  8.285 2.355 8.515 2.69 ;
      RECT  3.96 3.245 4.595 3.475 ;
      RECT  4.365 4.365 5.0 4.595 ;
      RECT  4.365 4.595 4.595 4.925 ;
      RECT  0.18 4.365 2.915 4.595 ;
      RECT  2.685 4.595 2.915 4.925 ;
      RECT  2.685 4.925 4.595 5.155 ;
  END
END MDN_AO311_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AO31_1
#      Description : One 3-input AND into 2-input OR
#      Equation    : X=(A1&A2&A3)|B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO31_1
  CLASS CORE ;
  FOREIGN MDN_AO31_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 4.365 4.06 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.905 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  0.0 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 5.715 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  4.66 3.245 5.715 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.67 1.005 2.76 1.235 ;
      RECT  3.19 1.565 4.04 1.795 ;
      RECT  3.81 1.795 4.04 2.405 ;
      RECT  3.81 2.405 5.21 2.635 ;
      RECT  3.81 2.635 4.04 3.245 ;
      RECT  3.81 3.245 4.3 3.475 ;
      RECT  3.245 4.365 3.475 4.925 ;
      RECT  0.905 4.925 3.475 5.155 ;
  END
END MDN_AO31_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AO31_2
#      Description : One 3-input AND into 2-input OR
#      Equation    : X=(A1&A2&A3)|B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO31_2
  CLASS CORE ;
  FOREIGN MDN_AO31_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 4.365 4.06 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  0.0 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 6.54 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  4.66 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  4.98 1.005 6.22 1.235 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  3.19 1.565 4.035 1.795 ;
      RECT  3.805 1.795 4.035 2.405 ;
      RECT  3.805 2.405 5.21 2.635 ;
      RECT  3.805 2.635 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
      RECT  3.245 4.365 3.475 4.925 ;
      RECT  0.95 4.925 3.475 5.155 ;
  END
END MDN_AO31_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AO31_4
#      Description : One 3-input AND into 2-input OR
#      Equation    : X=(A1&A2&A3)|B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO31_4
  CLASS CORE ;
  FOREIGN MDN_AO31_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 4.365 4.06 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  0.14 4.365 2.76 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  3.36 -0.14 4.035 0.14 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 8.78 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  4.66 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  1.67 1.005 2.76 1.235 ;
      RECT  3.19 1.565 4.03 1.795 ;
      RECT  3.8 1.795 4.03 2.405 ;
      RECT  3.8 2.405 6.33 2.635 ;
      RECT  3.8 2.635 4.03 3.245 ;
      RECT  3.8 3.245 4.3 3.475 ;
      RECT  7.11 2.405 8.565 2.635 ;
      RECT  3.245 4.365 3.475 4.925 ;
      RECT  0.95 4.925 3.475 5.155 ;
  END
END MDN_AO31_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AO32_1
#      Description : One 3-input AND one 2-input AND into 2-input OR
#      Equation    : X=(A1&A2&A3)|(B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO32_1
  CLASS CORE ;
  FOREIGN MDN_AO32_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 5.715 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.67 1.005 2.76 1.235 ;
      RECT  2.125 1.235 2.355 3.805 ;
      RECT  1.565 3.805 5.715 4.035 ;
      RECT  1.565 4.035 1.795 4.365 ;
      RECT  5.485 4.035 5.715 4.365 ;
      RECT  0.18 4.365 1.795 4.595 ;
      RECT  5.485 4.365 6.22 4.595 ;
      RECT  5.99 4.595 6.22 5.0 ;
      RECT  5.99 5.0 6.33 5.23 ;
      RECT  3.96 1.005 5.0 1.235 ;
      RECT  2.42 4.365 5.0 4.595 ;
      RECT  2.42 4.595 2.65 4.925 ;
      RECT  0.95 4.925 2.65 5.155 ;
  END
END MDN_AO32_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AO32_2
#      Description : One 3-input AND one 2-input AND into 2-input OR
#      Equation    : X=(A1&A2&A3)|(B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO32_2
  CLASS CORE ;
  FOREIGN MDN_AO32_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  4.925 -0.14 5.6 0.14 ;
      RECT  4.925 0.14 5.155 1.005 ;
      RECT  4.66 1.005 5.155 1.235 ;
      RECT  0.56 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 8.78 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  6.9 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 8.57 0.6 ;
      RECT  8.23 0.6 8.46 1.005 ;
      RECT  7.11 0.37 7.45 0.6 ;
      RECT  7.22 0.6 7.45 1.005 ;
      RECT  5.485 1.005 8.46 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  3.95 1.565 5.715 1.795 ;
      RECT  5.485 1.795 5.715 3.5 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  6.045 4.365 6.54 4.595 ;
      RECT  6.045 4.595 6.275 4.925 ;
      RECT  1.72 4.365 5.155 4.595 ;
      RECT  4.925 4.595 5.155 4.925 ;
      RECT  4.925 4.925 6.275 5.155 ;
  END
END MDN_AO32_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AO32_4
#      Description : One 3-input AND one 2-input AND into 2-input OR
#      Equation    : X=(A1&A2&A3)|(B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO32_4
  CLASS CORE ;
  FOREIGN MDN_AO32_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  7.28 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  4.925 -0.14 5.6 0.14 ;
      RECT  4.925 0.14 5.155 1.005 ;
      RECT  4.66 1.005 5.155 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 11.02 1.795 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  6.9 3.245 11.02 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  10.46 0.37 10.81 0.6 ;
      RECT  10.46 0.6 10.69 1.005 ;
      RECT  8.23 0.37 9.69 0.6 ;
      RECT  8.23 0.6 8.46 1.005 ;
      RECT  9.46 0.6 9.69 1.005 ;
      RECT  7.11 0.37 7.45 0.6 ;
      RECT  7.22 0.6 7.45 1.005 ;
      RECT  5.485 1.005 8.46 1.235 ;
      RECT  9.46 1.005 10.69 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  3.96 1.565 5.715 1.795 ;
      RECT  5.485 1.795 5.715 3.5 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  6.045 4.365 6.54 4.595 ;
      RECT  6.045 4.595 6.275 4.925 ;
      RECT  1.72 4.365 5.155 4.595 ;
      RECT  4.925 4.595 5.155 4.925 ;
      RECT  4.925 4.925 6.275 5.155 ;
  END
END MDN_AO32_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AO41_1
#      Description : One 4-input AND into 2-input OR
#      Equation    : X=(A1&A2&A3&A4)|B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO41_1
  CLASS CORE ;
  FOREIGN MDN_AO41_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A4
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  0.445 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  0.445 5.46 3.475 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  0.95 0.445 5.155 0.675 ;
      RECT  4.925 0.675 5.155 1.005 ;
      RECT  3.245 0.675 3.475 3.805 ;
      RECT  4.925 1.005 6.22 1.235 ;
      RECT  0.18 3.805 3.475 4.035 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  3.96 1.005 4.595 1.235 ;
      RECT  4.365 1.235 4.595 1.565 ;
      RECT  4.365 1.565 5.0 1.795 ;
      RECT  2.42 4.365 5.0 4.595 ;
      RECT  2.42 4.595 2.65 4.925 ;
      RECT  0.95 4.925 2.65 5.155 ;
  END
END MDN_AO41_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AO41_2
#      Description : One 4-input AND into 2-input OR
#      Equation    : X=(A1&A2&A3&A4)|B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO41_2
  CLASS CORE ;
  FOREIGN MDN_AO41_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A4
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.445 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  6.2 3.245 7.24 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.98 0.37 7.45 0.6 ;
      RECT  5.98 0.6 6.21 1.005 ;
      RECT  0.95 0.445 5.155 0.675 ;
      RECT  4.925 0.675 5.155 1.005 ;
      RECT  3.245 0.675 3.475 3.805 ;
      RECT  4.925 1.005 6.21 1.235 ;
      RECT  0.18 3.805 3.475 4.035 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  3.96 1.005 4.595 1.235 ;
      RECT  4.365 1.235 4.595 1.565 ;
      RECT  4.365 1.565 5.0 1.795 ;
      RECT  2.42 4.365 5.0 4.595 ;
      RECT  2.42 4.595 2.65 4.925 ;
      RECT  0.95 4.925 2.65 5.155 ;
  END
END MDN_AO41_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AO41_4
#      Description : One 4-input AND into 2-input OR
#      Equation    : X=(A1&A2&A3&A4)|B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AO41_4
  CLASS CORE ;
  FOREIGN MDN_AO41_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A4
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.445 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 9.48 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  6.2 3.245 9.48 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 9.69 0.6 ;
      RECT  8.23 0.6 8.46 1.005 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  7.215 0.6 7.445 1.005 ;
      RECT  0.95 0.445 5.155 0.675 ;
      RECT  4.925 0.675 5.155 1.005 ;
      RECT  3.245 0.675 3.475 3.805 ;
      RECT  4.925 1.005 6.22 1.235 ;
      RECT  7.215 1.005 8.46 1.235 ;
      RECT  0.18 3.805 3.475 4.035 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  3.96 1.005 4.595 1.235 ;
      RECT  4.365 1.235 4.595 1.565 ;
      RECT  4.365 1.565 5.0 1.795 ;
      RECT  2.42 4.365 5.0 4.595 ;
      RECT  2.42 4.595 2.65 4.925 ;
      RECT  0.95 4.925 2.65 5.155 ;
  END
END MDN_AO41_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AOAI211_1
#      Description : One 2-input AND into 2-input OR into 2-input NAND
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOAI211_1
  CLASS CORE ;
  FOREIGN MDN_AOAI211_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 4.65 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 1.565 ;
      RECT  1.005 1.565 2.76 1.795 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 1.005 4.3 1.235 ;
      RECT  3.245 1.235 3.475 3.53 ;
    END
    ANTENNADIFFAREA 2.086 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  2.125 0.445 3.53 0.675 ;
      RECT  2.125 0.675 2.355 1.005 ;
      RECT  1.72 1.005 2.355 1.235 ;
      RECT  0.18 4.365 2.76 4.595 ;
  END
END MDN_AOAI211_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AOAI211_2
#      Description : One 2-input AND into 2-input OR into 2-input NAND
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOAI211_2
  CLASS CORE ;
  FOREIGN MDN_AOAI211_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.605 1.565 8.01 1.795 ;
      RECT  6.605 1.795 6.835 4.365 ;
      RECT  4.66 4.365 8.78 4.595 ;
    END
    ANTENNADIFFAREA 4.686 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.83 0.445 3.53 0.675 ;
      RECT  1.83 0.675 2.06 1.005 ;
      RECT  0.18 1.005 2.06 1.235 ;
      RECT  2.42 1.005 8.78 1.235 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.07 4.595 4.3 4.925 ;
      RECT  4.065 4.925 5.77 5.155 ;
  END
END MDN_AOAI211_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AOAI211_3
#      Description : One 2-input AND into 2-input OR into 2-input NAND
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOAI211_3
  CLASS CORE ;
  FOREIGN MDN_AOAI211_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 6.3 2.355 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 9.66 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 2.125 13.02 2.355 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  10.525 4.365 11.02 4.595 ;
      RECT  10.525 4.595 10.755 5.46 ;
      RECT  10.08 5.46 10.755 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.88 -0.14 13.61 0.14 ;
      RECT  9.405 -0.14 10.08 0.14 ;
      RECT  9.405 0.14 9.635 1.005 ;
      RECT  9.14 1.005 9.635 1.235 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 2.76 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.525 1.565 12.49 1.795 ;
      RECT  10.525 1.795 10.755 3.805 ;
      RECT  9.965 3.805 11.875 4.035 ;
      RECT  11.645 4.035 11.875 4.365 ;
      RECT  9.965 4.035 10.195 4.925 ;
      RECT  11.645 4.365 13.26 4.595 ;
      RECT  7.67 4.925 10.195 5.155 ;
    END
    ANTENNADIFFAREA 6.448 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 11.93 0.6 ;
      RECT  0.95 0.445 5.77 0.675 ;
      RECT  9.965 1.005 13.26 1.235 ;
      RECT  9.965 1.235 10.195 1.565 ;
      RECT  3.96 1.005 8.515 1.235 ;
      RECT  8.285 1.235 8.515 1.565 ;
      RECT  8.285 1.565 10.195 1.795 ;
      RECT  0.18 4.365 9.48 4.595 ;
  END
END MDN_AOAI211_3
#-----------------------------------------------------------------------
#      Cell        : MDN_AOAI211_4
#      Description : One 2-input AND into 2-input OR into 2-input NAND
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOAI211_4
  CLASS CORE ;
  FOREIGN MDN_AOAI211_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  17.36 -0.14 18.09 0.14 ;
      RECT  11.76 -0.14 12.435 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.885 1.005 17.74 1.235 ;
      RECT  13.885 1.235 14.115 1.565 ;
      RECT  13.325 1.565 14.115 1.795 ;
      RECT  13.325 1.795 13.555 4.365 ;
      RECT  9.14 4.365 17.74 4.595 ;
    END
    ANTENNADIFFAREA 9.64 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  13.03 0.445 16.97 0.675 ;
      RECT  13.03 0.675 13.26 1.005 ;
      RECT  5.43 0.445 9.37 0.675 ;
      RECT  9.14 0.675 9.37 1.005 ;
      RECT  9.14 1.005 13.26 1.235 ;
      RECT  0.18 1.005 8.78 1.235 ;
      RECT  0.18 4.365 8.78 4.595 ;
      RECT  8.55 4.595 8.78 4.925 ;
      RECT  8.55 4.925 12.49 5.155 ;
  END
END MDN_AOAI211_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI211_1
#      Description : One 2-input AND into 3-input NOR
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI211_1
  CLASS CORE ;
  FOREIGN MDN_AOI211_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 4.365 4.06 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.695 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.72 1.005 4.3 1.235 ;
      RECT  3.805 1.235 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
    END
    ANTENNADIFFAREA 2.74 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 4.365 2.76 4.595 ;
  END
END MDN_AOI211_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI211_2
#      Description : One 2-input AND into 3-input NOR
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI211_2
  CLASS CORE ;
  FOREIGN MDN_AOI211_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  1.005 5.46 3.475 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  1.005 -0.14 2.41 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 8.78 1.235 ;
      RECT  6.605 1.235 6.835 3.245 ;
      RECT  6.605 3.245 8.01 3.475 ;
    END
    ANTENNADIFFAREA 5.156 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.815 0.445 3.53 0.675 ;
      RECT  1.815 0.675 2.045 1.005 ;
      RECT  0.18 1.005 2.06 1.235 ;
      RECT  0.18 4.365 6.54 4.595 ;
      RECT  8.285 4.365 8.78 4.595 ;
      RECT  8.285 4.595 8.515 4.925 ;
      RECT  6.955 4.34 7.185 4.925 ;
      RECT  5.43 4.925 8.515 5.155 ;
  END
END MDN_AOI211_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI211_3
#      Description : One 2-input AND into 3-input NOR
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI211_3
  CLASS CORE ;
  FOREIGN MDN_AOI211_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 7.42 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 16.38 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 11.9 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  17.36 5.46 18.09 5.74 ;
      RECT  7.165 4.925 8.01 5.155 ;
      RECT  7.165 5.155 7.395 5.46 ;
      RECT  5.43 4.925 6.275 5.155 ;
      RECT  6.045 5.155 6.275 5.46 ;
      RECT  6.045 5.46 7.395 5.74 ;
      RECT  2.685 4.925 3.53 5.155 ;
      RECT  2.685 5.155 2.915 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 2.915 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.005 16.2 1.235 ;
      RECT  13.325 1.235 13.555 3.245 ;
      RECT  13.325 3.245 16.2 3.475 ;
    END
    ANTENNADIFFAREA 8.22 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.805 0.445 8.01 0.675 ;
      RECT  3.805 0.675 4.035 1.005 ;
      RECT  0.18 1.005 4.035 1.235 ;
      RECT  0.18 4.365 8.515 4.595 ;
      RECT  8.285 4.595 8.515 4.925 ;
      RECT  8.285 4.925 12.49 5.155 ;
      RECT  9.14 4.365 12.995 4.595 ;
      RECT  12.765 4.595 12.995 4.925 ;
      RECT  12.765 4.925 16.97 5.155 ;
  END
END MDN_AOI211_3
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI211_4
#      Description : One 2-input AND into 3-input NOR
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI211_4
  CLASS CORE ;
  FOREIGN MDN_AOI211_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.685 ;
      RECT  9.38 2.685 13.02 2.915 ;
      RECT  10.5 2.125 10.78 2.685 ;
      RECT  11.62 2.125 11.9 2.685 ;
      RECT  12.74 2.125 13.02 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 9.13 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  11.76 -0.14 12.435 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.65 1.005 17.74 1.235 ;
      RECT  13.325 1.235 13.555 3.245 ;
      RECT  13.325 3.245 16.925 3.475 ;
    END
    ANTENNADIFFAREA 10.636 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  4.055 0.445 8.01 0.675 ;
      RECT  4.055 0.675 4.285 1.005 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  0.18 4.365 13.26 4.595 ;
      RECT  15.915 4.345 16.145 4.925 ;
      RECT  9.91 4.925 17.685 5.155 ;
      RECT  17.455 4.345 17.685 4.925 ;
  END
END MDN_AOI211_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI21_1
#      Description : One 2-input AND into 2-input NOR
#      Equation    : X=!((A1&A2)|B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI21_1
  CLASS CORE ;
  FOREIGN MDN_AOI21_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.525 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 3.53 ;
    END
    ANTENNADIFFAREA 2.7 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.14 4.365 2.76 4.595 ;
  END
END MDN_AOI21_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI21_2
#      Description : One 2-input AND into 2-input NOR
#      Equation    : X=!((A1&A2)|B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI21_2
  CLASS CORE ;
  FOREIGN MDN_AOI21_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  1.005 5.46 3.475 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  1.005 -0.14 2.41 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 6.54 1.235 ;
      RECT  4.365 1.235 4.595 3.245 ;
      RECT  4.365 3.245 5.77 3.475 ;
    END
    ANTENNADIFFAREA 3.928 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.83 0.445 3.53 0.675 ;
      RECT  1.83 0.675 2.06 1.005 ;
      RECT  0.17 1.005 2.06 1.235 ;
      RECT  0.14 4.365 5.005 4.595 ;
      RECT  4.775 4.595 5.005 4.925 ;
      RECT  4.775 4.925 6.485 5.155 ;
      RECT  6.255 4.34 6.485 4.925 ;
  END
END MDN_AOI21_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI21_3
#      Description : One 2-input AND into 2-input NOR
#      Equation    : X=!((A1&A2)|B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI21_3
  CLASS CORE ;
  FOREIGN MDN_AOI21_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 6.3 2.355 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 9.66 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 5.46 11.37 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  6.16 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  6.605 0.14 6.835 1.005 ;
      RECT  3.96 1.005 6.835 1.235 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.15 1.005 9.62 1.235 ;
      RECT  7.15 1.235 7.38 1.565 ;
      RECT  0.18 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  3.245 1.565 7.38 1.795 ;
      RECT  6.605 1.795 6.835 3.805 ;
      RECT  6.605 3.805 7.38 4.035 ;
      RECT  7.15 4.035 7.38 4.365 ;
      RECT  7.15 4.365 9.525 4.595 ;
    END
    ANTENNADIFFAREA 6.378 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 5.77 0.675 ;
      RECT  0.18 4.365 6.835 4.595 ;
      RECT  6.605 4.595 6.835 4.925 ;
      RECT  6.605 4.925 10.25 5.155 ;
  END
END MDN_AOI21_3
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI21_4
#      Description : One 2-input AND into 2-input NOR
#      Equation    : X=!((A1&A2)|B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI21_4
  CLASS CORE ;
  FOREIGN MDN_AOI21_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.88 5.46 13.61 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.695 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.64 1.005 13.26 1.235 ;
      RECT  8.845 1.235 9.075 3.245 ;
      RECT  8.845 3.245 12.49 3.475 ;
    END
    ANTENNADIFFAREA 8.18 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  4.07 0.445 8.01 0.675 ;
      RECT  4.07 0.675 4.3 1.005 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  0.14 4.365 13.26 4.595 ;
  END
END MDN_AOI21_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI21B_1
#      Description : One 2-input AND into 2-input NOR (other input inverted)
#      Equation    : X=!((A1&A2)|!B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI21B_1
  CLASS CORE ;
  FOREIGN MDN_AOI21B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.335 2.94 3.475 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 4.365 4.06 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.925 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.18 4.365 0.52 4.37 ;
      RECT  0.18 4.37 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 4.65 0.14 ;
      RECT  3.245 0.14 3.475 1.35 ;
      RECT  1.72 1.35 3.475 1.58 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 1.51 1.235 3.245 ;
      RECT  1.005 3.245 2.06 3.475 ;
    END
    ANTENNADIFFAREA 1.992 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.43 0.445 2.355 0.675 ;
      RECT  2.125 0.675 2.355 0.89 ;
      RECT  0.43 0.675 0.66 1.005 ;
      RECT  2.125 0.89 2.76 1.12 ;
      RECT  0.18 1.005 0.66 1.235 ;
      RECT  3.805 1.595 4.3 1.81 ;
      RECT  1.565 1.81 4.3 1.825 ;
      RECT  1.565 1.825 4.035 2.04 ;
      RECT  1.565 2.04 1.795 2.66 ;
      RECT  3.805 2.04 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
      RECT  2.125 4.365 2.76 4.595 ;
      RECT  2.125 4.595 2.355 4.955 ;
      RECT  0.95 4.955 2.355 5.185 ;
  END
END MDN_AOI21B_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI21B_2
#      Description : One 2-input AND into 2-input NOR (other input inverted)
#      Equation    : X=!((A1&A2)|!B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI21B_2
  CLASS CORE ;
  FOREIGN MDN_AOI21B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 4.365 7.42 5.0 ;
      RECT  7.11 5.0 7.45 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 4.595 1.235 ;
      RECT  4.365 1.235 4.595 1.565 ;
      RECT  4.365 1.565 6.54 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  4.365 3.245 6.58 3.475 ;
    END
    ANTENNADIFFAREA 4.252 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.83 0.445 3.53 0.675 ;
      RECT  1.83 0.675 2.06 1.005 ;
      RECT  0.18 1.005 2.06 1.235 ;
      RECT  6.955 1.565 7.185 2.41 ;
      RECT  4.87 2.41 7.185 2.64 ;
      RECT  6.955 2.64 7.185 3.485 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.07 4.595 4.3 4.925 ;
      RECT  4.07 4.925 5.77 5.155 ;
  END
END MDN_AOI21B_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI21B_3
#      Description : One 2-input AND into 2-input NOR (other input inverted)
#      Equation    : X=!((A1&A2)|!B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI21B_3
  CLASS CORE ;
  FOREIGN MDN_AOI21B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 7.42 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 4.06 2.355 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 5.46 11.37 5.74 ;
      RECT  6.9 4.365 7.395 4.595 ;
      RECT  7.165 4.595 7.395 5.46 ;
      RECT  6.72 5.46 7.395 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 -0.14 11.37 0.14 ;
      RECT  8.4 -0.14 9.52 0.14 ;
      RECT  8.845 0.14 9.075 1.005 ;
      RECT  8.44 1.005 10.25 1.235 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  5.43 0.445 7.955 0.675 ;
      RECT  7.725 0.675 7.955 1.565 ;
      RECT  7.72 1.565 11.02 1.795 ;
      RECT  9.965 1.795 10.195 3.805 ;
      RECT  8.44 3.805 10.195 4.035 ;
    END
    ANTENNADIFFAREA 5.786 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  9.35 0.37 10.805 0.6 ;
      RECT  1.72 1.005 7.24 1.235 ;
      RECT  8.23 2.405 9.69 2.635 ;
      RECT  8.23 2.635 8.46 3.245 ;
      RECT  5.485 3.245 8.46 3.475 ;
      RECT  5.485 3.475 5.715 3.805 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 3.805 ;
      RECT  1.005 3.805 5.715 4.035 ;
      RECT  1.005 4.035 1.235 4.365 ;
      RECT  0.18 4.365 1.235 4.595 ;
      RECT  6.31 3.805 7.86 4.035 ;
      RECT  6.31 4.035 6.54 4.365 ;
      RECT  7.63 4.035 7.86 4.365 ;
      RECT  1.72 4.365 6.54 4.595 ;
      RECT  7.63 4.365 11.02 4.595 ;
  END
END MDN_AOI21B_3
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI21B_4
#      Description : One 2-input AND into 2-input NOR (other input inverted)
#      Equation    : X=!((A1&A2)|!B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI21B_4
  CLASS CORE ;
  FOREIGN MDN_AOI21B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 4.365 14.14 5.0 ;
      RECT  13.83 5.0 14.17 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.905 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.83 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.695 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  12.205 0.14 12.435 0.695 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.005 11.315 1.235 ;
      RECT  11.085 1.235 11.315 1.565 ;
      RECT  11.085 1.565 13.26 1.795 ;
      RECT  11.085 1.795 11.315 3.245 ;
      RECT  9.14 3.245 13.26 3.475 ;
    END
    ANTENNADIFFAREA 8.504 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 11.93 0.6 ;
      RECT  4.07 0.445 8.01 0.675 ;
      RECT  4.07 0.675 4.3 1.005 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  13.58 1.565 13.96 1.795 ;
      RECT  13.58 1.795 13.81 2.405 ;
      RECT  11.59 2.405 13.81 2.635 ;
      RECT  13.58 2.635 13.81 3.245 ;
      RECT  13.58 3.245 13.96 3.475 ;
      RECT  9.34 2.405 10.595 2.635 ;
      RECT  0.18 4.365 9.075 4.595 ;
      RECT  8.845 4.595 9.075 4.925 ;
      RECT  8.845 4.925 12.49 5.155 ;
  END
END MDN_AOI21B_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI221_1
#      Description : Two 2-input ANDs into 3-input NOR
#      Equation    : X=!((A1&A2)|(B1&B2)|C)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI221_1
  CLASS CORE ;
  FOREIGN MDN_AOI221_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  2.24 -0.14 2.915 0.14 ;
      RECT  2.685 0.14 2.915 1.005 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.24 1.005 5.715 1.235 ;
      RECT  3.24 1.235 3.47 1.565 ;
      RECT  5.485 1.235 5.715 3.53 ;
      RECT  1.72 1.565 3.47 1.795 ;
    END
    ANTENNADIFFAREA 3.314 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.715 4.34 4.945 4.925 ;
      RECT  3.19 4.925 4.945 5.155 ;
  END
END MDN_AOI221_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI221_2
#      Description : Two 2-input ANDs into 3-input NOR
#      Equation    : X=!((A1&A2)|(B1&B2)|C)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI221_2
  CLASS CORE ;
  FOREIGN MDN_AOI221_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 10.78 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 5.46 11.37 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.165 1.005 11.02 1.235 ;
      RECT  7.165 1.235 7.395 1.565 ;
      RECT  8.845 1.235 9.075 3.245 ;
      RECT  2.42 1.005 4.035 1.235 ;
      RECT  3.805 1.235 4.035 1.565 ;
      RECT  3.805 1.565 7.395 1.795 ;
      RECT  8.845 3.245 10.25 3.475 ;
    END
    ANTENNADIFFAREA 5.156 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.83 0.445 3.53 0.675 ;
      RECT  1.83 0.675 2.06 1.005 ;
      RECT  0.175 1.005 2.06 1.235 ;
      RECT  6.605 0.445 8.01 0.675 ;
      RECT  6.605 0.675 6.835 1.005 ;
      RECT  4.66 1.005 6.835 1.235 ;
      RECT  0.18 4.365 8.78 4.595 ;
      RECT  9.195 4.35 9.425 4.925 ;
      RECT  5.43 4.925 10.965 5.155 ;
      RECT  10.735 4.35 10.965 4.925 ;
  END
END MDN_AOI221_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI221_4
#      Description : Two 2-input ANDs into 3-input NOR
#      Equation    : X=!((A1&A2)|(B1&B2)|C)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI221_4
  CLASS CORE ;
  FOREIGN MDN_AOI221_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.34 2.125 21.98 2.355 ;
      RECT  18.34 2.355 18.62 2.915 ;
      RECT  19.46 2.355 19.74 2.915 ;
      RECT  20.58 2.355 20.86 2.915 ;
      RECT  21.7 2.355 21.98 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.84 5.46 22.57 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 9.13 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.73 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.87 1.005 22.22 1.235 ;
      RECT  13.87 1.235 14.1 1.565 ;
      RECT  17.805 1.235 18.035 3.245 ;
      RECT  4.66 1.005 8.515 1.235 ;
      RECT  8.285 1.235 8.515 1.565 ;
      RECT  8.285 1.565 14.1 1.795 ;
      RECT  17.805 3.245 21.45 3.475 ;
    END
    ANTENNADIFFAREA 10.636 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  4.07 0.445 8.01 0.675 ;
      RECT  4.07 0.675 4.3 1.005 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  13.325 0.445 16.975 0.675 ;
      RECT  13.325 0.675 13.555 1.005 ;
      RECT  9.14 1.005 13.555 1.235 ;
      RECT  0.18 4.365 17.74 4.595 ;
      RECT  21.685 4.365 22.22 4.595 ;
      RECT  21.685 4.595 21.915 4.925 ;
      RECT  20.34 4.365 20.82 4.595 ;
      RECT  20.59 4.595 20.82 4.925 ;
      RECT  9.91 4.925 21.915 5.155 ;
  END
END MDN_AOI221_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI22_1
#      Description : Two 2-input ANDs into 2-input NOR
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI22_1
  CLASS CORE ;
  FOREIGN MDN_AOI22_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.865 1.235 5.46 ;
      RECT  1.005 5.46 2.41 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 -0.14 4.48 0.14 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 3.53 ;
    END
    ANTENNADIFFAREA 2.7 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.76 4.365 4.3 4.595 ;
      RECT  3.76 4.595 3.99 4.925 ;
      RECT  0.175 4.365 2.9 4.595 ;
      RECT  2.67 4.595 2.9 4.925 ;
      RECT  2.67 4.925 3.99 5.155 ;
  END
END MDN_AOI22_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI22_2
#      Description : Two 2-input ANDs into 2-input NOR
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI22_2
  CLASS CORE ;
  FOREIGN MDN_AOI22_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.865 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 6.27 1.235 ;
      RECT  6.04 1.235 6.27 1.565 ;
      RECT  6.04 1.565 6.835 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  5.43 3.245 8.01 3.475 ;
    END
    ANTENNADIFFAREA 5.4 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.83 0.445 3.53 0.675 ;
      RECT  1.83 0.675 2.06 1.005 ;
      RECT  0.18 1.005 2.06 1.235 ;
      RECT  5.43 0.445 6.835 0.675 ;
      RECT  6.605 0.675 6.835 1.005 ;
      RECT  6.605 1.005 8.78 1.235 ;
      RECT  8.245 4.365 8.78 4.595 ;
      RECT  8.245 4.595 8.475 4.925 ;
      RECT  6.005 4.365 7.38 4.595 ;
      RECT  6.005 4.595 6.235 4.925 ;
      RECT  7.15 4.595 7.38 4.925 ;
      RECT  0.18 4.365 5.14 4.375 ;
      RECT  0.18 4.375 5.155 4.595 ;
      RECT  4.925 4.595 5.155 4.925 ;
      RECT  4.925 4.925 6.235 5.155 ;
      RECT  7.15 4.925 8.475 5.155 ;
  END
END MDN_AOI22_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI22_3
#      Description : Two 2-input ANDs into 2-input NOR
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI22_3
  CLASS CORE ;
  FOREIGN MDN_AOI22_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 9.66 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 13.02 2.355 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 6.3 2.355 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.88 5.46 13.61 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.32 -0.14 13.61 0.14 ;
      RECT  12.765 0.14 12.995 1.005 ;
      RECT  10.66 1.005 13.26 1.235 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 2.76 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.96 1.005 9.48 1.235 ;
      RECT  6.605 1.235 6.835 3.805 ;
      RECT  6.605 3.805 7.395 4.035 ;
      RECT  7.165 4.035 7.395 4.365 ;
      RECT  7.165 4.365 13.26 4.595 ;
    END
    ANTENNADIFFAREA 9.072 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.92 0.445 5.77 0.675 ;
      RECT  7.67 0.445 12.49 0.675 ;
      RECT  0.18 4.365 6.835 4.595 ;
      RECT  6.605 4.595 6.835 4.925 ;
      RECT  6.605 4.925 12.49 5.155 ;
  END
END MDN_AOI22_3
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI22_4
#      Description : Two 2-input ANDs into 2-input NOR
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI22_4
  CLASS CORE ;
  FOREIGN MDN_AOI22_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  17.36 5.46 18.09 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.65 1.005 12.995 1.235 ;
      RECT  12.765 1.235 12.995 1.565 ;
      RECT  12.765 1.565 13.555 1.795 ;
      RECT  13.325 1.795 13.555 4.365 ;
      RECT  9.14 4.365 17.74 4.595 ;
    END
    ANTENNADIFFAREA 12.096 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  4.07 0.445 8.01 0.675 ;
      RECT  4.07 0.675 4.3 1.005 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  9.895 0.445 13.555 0.675 ;
      RECT  13.325 0.675 13.555 1.005 ;
      RECT  13.325 1.005 17.74 1.235 ;
      RECT  0.18 4.365 8.78 4.595 ;
      RECT  8.55 4.595 8.78 4.925 ;
      RECT  8.55 4.925 16.97 5.155 ;
  END
END MDN_AOI22_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI311_1
#      Description : One 3-input AND into 3-input NOR
#      Equation    : X=!((A1&A2&A3)|B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI311_1
  CLASS CORE ;
  FOREIGN MDN_AOI311_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 4.365 6.3 5.0 ;
      RECT  5.99 5.0 6.33 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  1.005 5.46 3.475 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  1.005 -0.14 2.41 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.96 1.005 6.54 1.235 ;
      RECT  6.045 1.235 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 2.74 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.67 1.005 2.76 1.235 ;
      RECT  1.72 4.365 5.0 4.595 ;
  END
END MDN_AOI311_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI311_2
#      Description : One 3-input AND into 3-input NOR
#      Equation    : X=!((A1&A2&A3)|B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI311_2
  CLASS CORE ;
  FOREIGN MDN_AOI311_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 10.78 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 5.46 11.37 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.615 1.005 11.02 1.235 ;
      RECT  8.845 1.235 9.075 3.245 ;
      RECT  8.845 3.245 10.25 3.475 ;
    END
    ANTENNADIFFAREA 5.156 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.445 5.77 0.675 ;
      RECT  0.14 1.005 4.3 1.235 ;
      RECT  0.18 4.365 8.78 4.595 ;
      RECT  10.525 4.365 11.02 4.595 ;
      RECT  10.525 4.595 10.755 4.925 ;
      RECT  9.195 4.34 9.425 4.925 ;
      RECT  7.63 4.925 10.755 5.155 ;
  END
END MDN_AOI311_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI311_4
#      Description : One 3-input AND into 3-input NOR
#      Equation    : X=!((A1&A2&A3)|B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI311_4
  CLASS CORE ;
  FOREIGN MDN_AOI311_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.34 2.125 21.98 2.355 ;
      RECT  18.34 2.355 18.62 2.915 ;
      RECT  19.46 2.355 19.74 2.915 ;
      RECT  20.58 2.355 20.86 2.915 ;
      RECT  21.7 2.355 21.98 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.84 5.46 22.57 5.74 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.695 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  14.445 -0.14 16.915 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.14 1.005 22.22 1.235 ;
      RECT  17.805 1.235 18.035 3.245 ;
      RECT  17.805 3.245 21.45 3.475 ;
    END
    ANTENNADIFFAREA 10.636 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.445 12.49 0.675 ;
      RECT  0.14 1.005 8.78 1.235 ;
      RECT  0.18 4.365 17.74 4.595 ;
      RECT  20.045 4.365 22.22 4.595 ;
      RECT  20.045 4.595 20.275 4.925 ;
      RECT  14.39 4.925 20.275 5.155 ;
  END
END MDN_AOI311_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI31_1
#      Description : One 3-input AND into 2-input NOR
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI31_1
  CLASS CORE ;
  FOREIGN MDN_AOI31_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  0.14 4.365 2.76 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 -0.14 4.48 0.14 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 1.51 3.475 3.245 ;
      RECT  3.245 3.245 4.3 3.475 ;
    END
    ANTENNADIFFAREA 1.992 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  0.95 4.925 3.53 5.155 ;
  END
END MDN_AOI31_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI31_2
#      Description : One 3-input AND into 2-input NOR
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI31_2
  CLASS CORE ;
  FOREIGN MDN_AOI31_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  1.005 5.46 3.475 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.62 1.005 8.78 1.235 ;
      RECT  6.605 1.235 6.835 3.245 ;
      RECT  6.605 3.245 8.01 3.475 ;
    END
    ANTENNADIFFAREA 3.928 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.145 0.445 5.77 0.675 ;
      RECT  0.13 1.005 4.3 1.235 ;
      RECT  0.13 4.365 7.24 4.595 ;
      RECT  7.01 4.595 7.24 4.925 ;
      RECT  7.01 4.925 8.725 5.155 ;
      RECT  8.495 4.34 8.725 4.925 ;
  END
END MDN_AOI31_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI31_3
#      Description : One 3-input AND into 2-input NOR
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI31_3
  CLASS CORE ;
  FOREIGN MDN_AOI31_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 9.66 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 6.3 2.355 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 13.02 2.355 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.88 5.46 13.61 5.74 ;
      RECT  9.195 4.31 9.425 5.46 ;
      RECT  8.96 5.46 9.52 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.32 -0.14 13.61 0.14 ;
      RECT  12.765 0.14 12.995 1.005 ;
      RECT  10.66 1.005 13.26 1.235 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 2.76 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.67 0.445 12.49 0.675 ;
      RECT  9.965 0.675 10.195 3.245 ;
      RECT  9.965 3.245 10.755 3.475 ;
      RECT  10.525 3.475 10.755 4.365 ;
      RECT  10.525 4.365 13.26 4.595 ;
    END
    ANTENNADIFFAREA 5.976 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.92 0.445 5.77 0.675 ;
      RECT  3.96 1.005 9.48 1.235 ;
      RECT  8.285 3.805 10.195 4.035 ;
      RECT  8.285 4.035 8.515 4.365 ;
      RECT  9.965 4.035 10.195 4.925 ;
      RECT  0.18 4.365 8.515 4.595 ;
      RECT  9.965 4.925 12.49 5.155 ;
  END
END MDN_AOI31_3
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI31_4
#      Description : One 3-input AND into 2-input NOR
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI31_4
  CLASS CORE ;
  FOREIGN MDN_AOI31_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  17.36 5.46 18.09 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.13 1.005 17.74 1.235 ;
      RECT  13.325 1.235 13.555 3.245 ;
      RECT  13.325 3.245 16.97 3.475 ;
    END
    ANTENNADIFFAREA 8.18 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.445 12.49 0.675 ;
      RECT  0.14 1.005 8.78 1.235 ;
      RECT  0.14 4.365 13.555 4.595 ;
      RECT  13.325 4.595 13.555 4.925 ;
      RECT  13.325 4.925 17.685 5.155 ;
      RECT  15.915 4.34 16.145 4.925 ;
      RECT  17.455 4.34 17.685 4.925 ;
  END
END MDN_AOI31_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI32_1
#      Description : One 3-input AND one 2-input AND into into 2-input NOR
#      Equation    : X=!((A1&A2&A3)|(B1&B2))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI32_1
  CLASS CORE ;
  FOREIGN MDN_AOI32_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  1.005 5.46 3.475 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 -0.14 6.89 0.14 ;
      RECT  6.045 0.14 6.275 1.005 ;
      RECT  6.045 1.005 6.54 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.19 0.445 4.595 0.675 ;
      RECT  4.365 0.675 4.595 1.005 ;
      RECT  4.365 1.005 5.715 1.235 ;
      RECT  5.485 1.235 5.715 3.53 ;
    END
    ANTENNADIFFAREA 3.18 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  0.18 4.365 6.54 4.595 ;
  END
END MDN_AOI32_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI32_2
#      Description : One 3-input AND one 2-input AND into into 2-input NOR
#      Equation    : X=!((A1&A2&A3)|(B1&B2))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI32_2
  CLASS CORE ;
  FOREIGN MDN_AOI32_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 10.78 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 5.46 11.37 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.005 8.78 1.235 ;
      RECT  6.605 1.235 6.835 3.805 ;
      RECT  6.605 3.805 7.09 4.035 ;
      RECT  6.86 4.035 7.09 4.365 ;
      RECT  6.86 4.365 11.02 4.595 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.445 5.77 0.675 ;
      RECT  7.67 0.445 9.37 0.675 ;
      RECT  9.14 0.675 9.37 1.005 ;
      RECT  9.14 1.005 11.02 1.235 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  0.18 4.365 6.54 4.595 ;
      RECT  6.31 4.595 6.54 4.925 ;
      RECT  6.31 4.925 10.25 5.155 ;
  END
END MDN_AOI32_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI32_4
#      Description : One 3-input AND one 2-input AND into into 2-input NOR
#      Equation    : X=!((A1&A2&A3)|(B1&B2))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI32_4
  CLASS CORE ;
  FOREIGN MDN_AOI32_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.34 2.125 21.98 2.355 ;
      RECT  18.34 2.355 18.62 2.915 ;
      RECT  19.46 2.355 19.74 2.915 ;
      RECT  20.58 2.355 20.86 2.915 ;
      RECT  21.7 2.355 21.98 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.84 5.46 22.57 5.74 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.73 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  10.64 -0.14 11.76 0.14 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.13 1.005 17.74 1.235 ;
      RECT  13.325 1.235 13.555 3.805 ;
      RECT  13.325 3.805 14.1 4.035 ;
      RECT  13.87 4.035 14.1 4.365 ;
      RECT  13.87 4.365 22.22 4.595 ;
    END
    ANTENNADIFFAREA 12.096 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.445 12.49 0.675 ;
      RECT  14.39 0.445 18.33 0.675 ;
      RECT  18.1 0.675 18.33 1.005 ;
      RECT  18.1 1.005 22.22 1.235 ;
      RECT  0.18 1.005 8.78 1.235 ;
      RECT  0.18 4.365 13.555 4.595 ;
      RECT  13.325 4.595 13.555 4.925 ;
      RECT  13.325 4.925 21.45 5.155 ;
  END
END MDN_AOI32_4
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI41_1
#      Description : One 4-input AND into 2-input NOR
#      Equation    : X=!((A1&A2&A3&A4)|B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI41_1
  CLASS CORE ;
  FOREIGN MDN_AOI41_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A4
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  1.005 5.46 3.475 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.96 1.005 4.3 1.01 ;
      RECT  3.96 1.01 5.715 1.24 ;
      RECT  4.66 1.005 5.0 1.01 ;
      RECT  5.485 1.005 5.715 1.01 ;
      RECT  5.485 1.24 5.715 3.53 ;
    END
    ANTENNADIFFAREA 2.7 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  0.18 4.365 5.0 4.595 ;
  END
END MDN_AOI41_1
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI41_2
#      Description : One 4-input AND into 2-input NOR
#      Equation    : X=!((A1&A2&A3&A4)|B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI41_2
  CLASS CORE ;
  FOREIGN MDN_AOI41_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.115 8.54 2.345 ;
      RECT  7.14 2.345 7.42 2.915 ;
      RECT  8.26 2.345 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.115 6.3 2.345 ;
      RECT  4.9 2.345 5.18 2.915 ;
      RECT  6.02 2.345 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.115 4.06 2.345 ;
      RECT  2.66 2.345 2.94 2.915 ;
      RECT  3.78 2.345 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.115 1.82 2.345 ;
      RECT  0.42 2.345 0.7 2.915 ;
      RECT  1.54 2.345 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A4
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.115 10.78 2.345 ;
      RECT  9.38 2.345 9.66 2.915 ;
      RECT  10.5 2.345 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 5.46 11.37 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.855 1.005 11.02 1.235 ;
      RECT  8.845 1.235 9.075 3.245 ;
      RECT  8.845 3.245 10.25 3.475 ;
    END
    ANTENNADIFFAREA 3.928 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.445 4.85 0.675 ;
      RECT  4.62 0.675 4.85 1.005 ;
      RECT  4.62 1.005 6.54 1.235 ;
      RECT  5.43 0.445 8.01 0.675 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  0.14 4.365 9.62 4.595 ;
      RECT  9.39 4.595 9.62 4.925 ;
      RECT  9.39 4.925 10.965 5.155 ;
      RECT  10.735 4.34 10.965 4.925 ;
  END
END MDN_AOI41_2
#-----------------------------------------------------------------------
#      Cell        : MDN_AOI41_4
#      Description : One 4-input AND into 2-input NOR
#      Equation    : X=!((A1&A2&A3&A4)|B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_AOI41_4
  CLASS CORE ;
  FOREIGN MDN_AOI41_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A4
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.34 2.125 21.98 2.355 ;
      RECT  18.34 2.355 18.62 2.915 ;
      RECT  19.46 2.355 19.74 2.915 ;
      RECT  20.58 2.355 20.86 2.915 ;
      RECT  21.7 2.355 21.98 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.84 5.46 22.57 5.74 ;
      RECT  14.445 4.87 14.675 5.46 ;
      RECT  14.445 5.46 16.915 5.74 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.695 ;
      RECT  18.925 -0.14 19.6 0.14 ;
      RECT  18.925 0.14 19.155 0.695 ;
      RECT  10.64 -0.14 11.76 0.14 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.61 1.005 22.22 1.235 ;
      RECT  17.805 1.235 18.035 3.245 ;
      RECT  17.805 3.245 21.45 3.475 ;
    END
    ANTENNADIFFAREA 8.18 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.445 12.49 0.675 ;
      RECT  13.03 0.445 16.97 0.675 ;
      RECT  13.03 0.675 13.26 1.005 ;
      RECT  9.14 1.005 13.26 1.235 ;
      RECT  0.18 1.005 8.78 1.235 ;
      RECT  21.685 4.365 22.22 4.595 ;
      RECT  21.685 4.595 21.915 4.925 ;
      RECT  20.34 4.365 20.82 4.595 ;
      RECT  20.59 4.595 20.82 4.925 ;
      RECT  0.18 4.365 18.035 4.595 ;
      RECT  17.805 4.595 18.035 4.925 ;
      RECT  17.805 4.925 21.915 5.155 ;
  END
END MDN_AOI41_4
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_1
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_1
  CLASS CORE ;
  FOREIGN MDN_BUF_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.24 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 4.365 0.7 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 2.24 5.74 ;
      LAYER VIA12 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 2.24 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 1.74 1.235 ;
      RECT  0.44 1.235 0.67 3.245 ;
      RECT  0.18 3.245 0.67 3.475 ;
  END
END MDN_BUF_1
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_12
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_12
  CLASS CORE ;
  FOREIGN MDN_BUF_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.92 1.4 16.52 1.96 ;
      RECT  15.96 1.96 16.52 3.08 ;
      RECT  3.96 3.08 16.52 3.64 ;
    END
    ANTENNADIFFAREA 18.144 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  14.95 0.37 16.41 0.6 ;
      RECT  0.18 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 2.405 ;
      RECT  3.245 2.405 15.29 2.635 ;
      RECT  3.245 2.635 3.475 3.805 ;
      RECT  0.18 3.805 3.475 4.035 ;
  END
END MDN_BUF_12
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_16
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_16
  CLASS CORE ;
  FOREIGN MDN_BUF_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 2.94 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
      RECT  2.66 2.125 2.94 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.905 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.905 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  16.685 4.905 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  14.445 4.905 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  9.965 4.905 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.905 12.435 5.46 ;
      RECT  7.725 4.905 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.905 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.905 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.905 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.695 ;
      RECT  18.925 -0.14 19.6 0.14 ;
      RECT  18.925 0.14 19.155 0.695 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.695 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.695 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 22.22 1.795 ;
      RECT  20.045 1.795 20.275 3.245 ;
      RECT  4.66 3.245 22.22 3.475 ;
    END
    ANTENNADIFFAREA 24.192 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.09 0.375 ;
      RECT  3.74 0.375 4.09 0.6 ;
      RECT  3.74 0.6 3.97 1.005 ;
      RECT  2.63 0.37 2.99 0.6 ;
      RECT  2.76 0.6 2.99 1.005 ;
      RECT  2.76 1.005 3.97 1.235 ;
      RECT  19.43 0.37 20.89 0.6 ;
      RECT  0.18 1.005 2.355 1.235 ;
      RECT  2.125 1.235 2.355 1.565 ;
      RECT  2.125 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 2.405 ;
      RECT  3.805 2.405 19.77 2.635 ;
      RECT  3.805 2.635 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
      RECT  3.805 3.475 4.035 3.805 ;
      RECT  0.18 3.805 4.035 4.035 ;
      RECT  20.55 2.405 22.01 2.635 ;
  END
END MDN_BUF_16
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_2
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_2
  CLASS CORE ;
  FOREIGN MDN_BUF_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 4.365 0.7 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 4.65 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  1.005 5.46 1.68 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.72 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 3.245 ;
      RECT  1.72 3.245 3.475 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.565 0.675 1.795 ;
      RECT  0.445 1.795 0.675 2.125 ;
      RECT  0.445 2.125 2.915 2.355 ;
      RECT  1.565 2.355 1.795 2.69 ;
      RECT  2.685 2.355 2.915 2.69 ;
      RECT  0.445 2.355 0.675 3.245 ;
      RECT  0.18 3.245 0.675 3.475 ;
  END
END MDN_BUF_2
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_24
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_24
  CLASS CORE ;
  FOREIGN MDN_BUF_24 0 0 ;
  ORIGIN 0 0 ;
  SIZE 33.6 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 5.18 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  32.365 4.87 32.595 5.46 ;
      RECT  32.365 5.46 33.77 5.74 ;
      RECT  30.125 4.9 30.355 5.46 ;
      RECT  29.68 5.46 30.355 5.74 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.645 5.46 28.115 5.74 ;
      RECT  27.885 4.9 28.115 5.46 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  22.96 5.46 23.635 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  20.72 5.46 21.395 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 19.155 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 33.6 5.74 ;
      LAYER VIA12 ;
      RECT  32.63 5.47 32.89 5.73 ;
      RECT  33.19 5.47 33.45 5.73 ;
      RECT  29.83 5.47 30.09 5.73 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  27.03 5.47 27.29 5.73 ;
      RECT  27.59 5.47 27.85 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  18.07 5.47 18.33 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  32.365 -0.14 33.77 0.14 ;
      RECT  32.365 0.14 32.595 0.715 ;
      RECT  29.68 -0.14 30.355 0.14 ;
      RECT  30.125 0.14 30.355 0.715 ;
      RECT  25.645 -0.14 28.115 0.14 ;
      RECT  25.645 0.14 25.875 0.715 ;
      RECT  27.885 0.14 28.115 0.715 ;
      RECT  22.96 -0.14 23.635 0.14 ;
      RECT  23.405 0.14 23.635 0.715 ;
      RECT  20.72 -0.14 21.395 0.14 ;
      RECT  21.165 0.14 21.395 0.715 ;
      RECT  16.685 -0.14 19.155 0.14 ;
      RECT  16.685 0.14 16.915 0.715 ;
      RECT  18.925 0.14 19.155 0.715 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.715 ;
      RECT  11.76 -0.14 12.435 0.14 ;
      RECT  12.205 0.14 12.435 0.715 ;
      RECT  7.725 -0.14 10.195 0.14 ;
      RECT  7.725 0.14 7.955 0.715 ;
      RECT  9.965 0.14 10.195 0.715 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 33.6 0.14 ;
      LAYER VIA12 ;
      RECT  32.63 -0.13 32.89 0.13 ;
      RECT  33.19 -0.13 33.45 0.13 ;
      RECT  29.83 -0.13 30.09 0.13 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  27.03 -0.13 27.29 0.13 ;
      RECT  27.59 -0.13 27.85 0.13 ;
      RECT  23.11 -0.13 23.37 0.13 ;
      RECT  20.87 -0.13 21.13 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  18.07 -0.13 18.33 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.955 0.945 32.11 1.51 ;
      RECT  6.955 1.51 33.365 1.85 ;
      RECT  6.955 1.85 32.11 2.055 ;
      RECT  31.0 2.055 32.11 2.98 ;
      RECT  6.955 2.98 32.11 3.19 ;
      RECT  6.955 3.19 33.365 3.53 ;
      RECT  6.955 3.53 32.11 3.92 ;
      RECT  6.955 3.92 32.105 4.09 ;
    END
    ANTENNADIFFAREA 36.288 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  4.87 0.37 5.23 0.6 ;
      RECT  5.0 0.6 5.23 1.005 ;
      RECT  5.0 1.005 6.22 1.235 ;
      RECT  0.17 1.005 4.595 1.235 ;
      RECT  4.365 1.235 4.595 1.565 ;
      RECT  4.365 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 2.405 ;
      RECT  6.045 2.405 30.77 2.635 ;
      RECT  6.045 2.635 6.275 3.805 ;
      RECT  0.17 3.805 6.54 4.035 ;
      RECT  31.88 4.365 33.09 4.595 ;
      RECT  31.88 4.595 32.11 5.0 ;
      RECT  32.86 4.595 33.09 5.0 ;
      RECT  30.63 5.0 32.11 5.23 ;
      RECT  32.86 5.0 33.21 5.23 ;
  END
END MDN_BUF_24
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_3
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_3
  CLASS CORE ;
  FOREIGN MDN_BUF_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 4.365 0.7 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 4.65 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  1.005 5.46 1.68 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      RECT  3.245 0.14 3.475 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.72 1.565 4.3 1.795 ;
      RECT  2.125 1.795 2.355 3.245 ;
      RECT  1.72 3.245 4.3 3.475 ;
    END
    ANTENNADIFFAREA 4.536 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 2.99 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 1.74 1.235 ;
      RECT  0.445 1.235 0.675 3.245 ;
      RECT  0.18 3.245 0.675 3.475 ;
      RECT  2.685 2.125 4.035 2.355 ;
      RECT  2.685 2.355 2.915 2.69 ;
      RECT  3.805 2.355 4.035 2.69 ;
  END
END MDN_BUF_3
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_4
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_4
  CLASS CORE ;
  FOREIGN MDN_BUF_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  1.005 -0.14 1.68 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 6.54 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  2.42 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.75 0.37 5.23 0.6 ;
      RECT  5.0 0.6 5.23 1.005 ;
      RECT  5.0 1.005 6.22 1.235 ;
      RECT  1.525 1.565 2.06 1.795 ;
      RECT  1.525 1.795 1.755 2.405 ;
      RECT  1.525 2.405 4.09 2.635 ;
      RECT  1.525 2.635 1.755 3.245 ;
      RECT  1.525 3.245 2.06 3.475 ;
  END
END MDN_BUF_4
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_6
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_6
  CLASS CORE ;
  FOREIGN MDN_BUF_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 9.13 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  2.685 1.235 2.915 1.565 ;
      RECT  2.685 1.565 8.78 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  2.685 3.245 8.78 3.475 ;
      RECT  2.685 3.475 2.915 4.365 ;
      RECT  2.42 4.365 2.915 4.595 ;
    END
    ANTENNADIFFAREA 9.072 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 2.125 ;
      RECT  2.125 2.125 6.275 2.355 ;
      RECT  2.685 2.355 2.915 2.69 ;
      RECT  3.805 2.355 4.035 2.69 ;
      RECT  4.925 2.355 5.155 2.69 ;
      RECT  6.045 2.355 6.275 2.69 ;
      RECT  2.125 2.355 2.355 3.805 ;
      RECT  1.565 3.805 2.355 4.035 ;
      RECT  1.565 4.035 1.795 4.365 ;
      RECT  0.18 4.365 1.795 4.595 ;
      RECT  7.165 2.125 8.515 2.355 ;
      RECT  7.165 2.355 7.395 2.69 ;
      RECT  8.285 2.355 8.515 2.69 ;
  END
END MDN_BUF_6
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_8
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_8
  CLASS CORE ;
  FOREIGN MDN_BUF_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  2.685 1.235 2.915 1.565 ;
      RECT  2.685 1.565 11.02 1.795 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  2.685 3.245 11.02 3.475 ;
      RECT  2.685 3.475 2.915 4.365 ;
      RECT  2.42 4.365 2.915 4.595 ;
    END
    ANTENNADIFFAREA 12.096 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 9.69 0.6 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 2.125 ;
      RECT  2.125 2.125 8.515 2.355 ;
      RECT  2.685 2.355 2.915 2.69 ;
      RECT  3.805 2.355 4.035 2.69 ;
      RECT  4.925 2.355 5.155 2.69 ;
      RECT  6.045 2.355 6.275 2.69 ;
      RECT  7.165 2.355 7.395 2.69 ;
      RECT  8.285 2.355 8.515 2.69 ;
      RECT  2.125 2.355 2.355 3.805 ;
      RECT  1.565 3.805 2.355 4.035 ;
      RECT  1.565 4.035 1.795 4.365 ;
      RECT  0.18 4.365 1.795 4.595 ;
      RECT  9.405 2.125 10.755 2.355 ;
      RECT  9.405 2.355 9.635 2.69 ;
      RECT  10.525 2.355 10.755 2.69 ;
  END
END MDN_BUF_8
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_AS_1
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_AS_1
  CLASS CORE ;
  FOREIGN MDN_BUF_AS_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 1.565 2.06 1.795 ;
      RECT  1.54 1.795 1.795 2.125 ;
      RECT  1.54 2.125 4.06 2.355 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNADIFFAREA 0.614 ;
    ANTENNAGATEAREA 1.701 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 5.715 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.695 ;
      RECT  5.485 0.14 5.715 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 1.565 6.545 1.795 ;
      RECT  5.485 1.795 5.715 3.805 ;
      RECT  4.66 3.805 6.54 4.035 ;
    END
    ANTENNADIFFAREA 2.41 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.955 1.565 4.595 1.795 ;
      RECT  4.365 1.795 4.595 2.405 ;
      RECT  4.365 2.405 5.21 2.635 ;
      RECT  4.365 2.635 4.595 3.245 ;
      RECT  2.38 3.245 4.595 3.475 ;
      RECT  5.0 4.365 6.22 4.595 ;
      RECT  5.0 4.595 5.23 5.0 ;
      RECT  5.99 4.595 6.22 5.0 ;
      RECT  4.87 5.0 5.23 5.23 ;
      RECT  5.99 5.0 6.33 5.23 ;
  END
END MDN_BUF_AS_1
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_AS_12
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_AS_12
  CLASS CORE ;
  FOREIGN MDN_BUF_AS_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 33.6 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.125 ;
      RECT  0.42 2.125 6.275 2.355 ;
      RECT  6.045 2.355 6.275 2.69 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
    END
    ANTENNADIFFAREA 0.614 ;
    ANTENNAGATEAREA 3.402 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  32.925 4.365 33.42 4.595 ;
      RECT  32.925 4.595 33.155 5.46 ;
      RECT  32.925 5.46 33.77 5.74 ;
      RECT  31.54 4.365 32.035 4.595 ;
      RECT  31.805 4.595 32.035 5.46 ;
      RECT  31.19 5.46 32.035 5.74 ;
      RECT  27.885 4.9 28.115 5.46 ;
      RECT  27.885 5.46 30.355 5.74 ;
      RECT  30.125 4.9 30.355 5.46 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.645 5.46 26.32 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 23.635 5.74 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 16.915 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 33.6 5.74 ;
      LAYER VIA12 ;
      RECT  33.19 5.47 33.45 5.73 ;
      RECT  31.51 5.47 31.77 5.73 ;
      RECT  28.15 5.47 28.41 5.73 ;
      RECT  28.71 5.47 28.97 5.73 ;
      RECT  29.27 5.47 29.53 5.73 ;
      RECT  29.83 5.47 30.09 5.73 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  22.55 5.47 22.81 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  30.125 -0.14 33.77 0.14 ;
      RECT  30.125 0.14 30.355 0.7 ;
      RECT  27.885 -0.14 28.56 0.14 ;
      RECT  27.885 0.14 28.115 0.7 ;
      RECT  23.405 -0.14 25.875 0.14 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  25.645 0.14 25.875 0.7 ;
      RECT  20.72 -0.14 21.395 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  12.88 -0.14 14.0 0.14 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 33.6 0.14 ;
      LAYER VIA12 ;
      RECT  30.39 -0.13 30.65 0.13 ;
      RECT  30.95 -0.13 31.21 0.13 ;
      RECT  31.51 -0.13 31.77 0.13 ;
      RECT  32.07 -0.13 32.33 0.13 ;
      RECT  32.63 -0.13 32.89 0.13 ;
      RECT  33.19 -0.13 33.45 0.13 ;
      RECT  28.15 -0.13 28.41 0.13 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  24.79 -0.13 25.05 0.13 ;
      RECT  25.35 -0.13 25.61 0.13 ;
      RECT  20.87 -0.13 21.13 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  16.565 1.49 32.155 1.96 ;
      RECT  16.565 1.96 17.035 3.08 ;
      RECT  31.685 1.96 32.155 3.08 ;
      RECT  8.32 3.08 32.65 3.085 ;
      RECT  8.165 3.085 32.65 3.55 ;
      RECT  8.165 3.55 8.635 3.64 ;
      RECT  6.955 3.64 8.635 4.11 ;
    END
    ANTENNADIFFAREA 28.596 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  16.07 0.37 18.65 0.6 ;
      RECT  30.63 0.37 33.21 0.6 ;
      RECT  3.94 1.565 6.835 1.795 ;
      RECT  6.605 1.795 6.835 2.405 ;
      RECT  6.605 2.405 16.225 2.635 ;
      RECT  6.605 2.635 6.835 3.21 ;
      RECT  6.005 3.21 6.835 3.44 ;
      RECT  6.005 3.44 6.235 3.805 ;
      RECT  0.17 3.805 6.235 4.035 ;
      RECT  17.385 2.405 30.97 2.635 ;
  END
END MDN_BUF_AS_12
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_AS_16
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_AS_16
  CLASS CORE ;
  FOREIGN MDN_BUF_AS_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 44.8 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.125 ;
      RECT  0.42 2.125 6.3 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNADIFFAREA 0.614 ;
    ANTENNAGATEAREA 4.536 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  43.565 4.9 43.795 5.46 ;
      RECT  43.565 5.46 44.97 5.74 ;
      RECT  41.325 4.9 41.555 5.46 ;
      RECT  41.325 5.46 42.0 5.74 ;
      RECT  39.085 4.9 39.315 5.46 ;
      RECT  38.64 5.46 39.315 5.74 ;
      RECT  36.845 4.9 37.075 5.46 ;
      RECT  36.845 5.46 37.52 5.74 ;
      RECT  34.605 4.9 34.835 5.46 ;
      RECT  34.16 5.46 34.835 5.74 ;
      RECT  32.365 4.9 32.595 5.46 ;
      RECT  32.365 5.46 33.04 5.74 ;
      RECT  27.885 4.9 28.115 5.46 ;
      RECT  27.885 5.46 30.355 5.74 ;
      RECT  30.125 4.9 30.355 5.46 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.2 5.46 25.875 5.74 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.08 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  20.72 5.46 21.395 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 16.915 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 5.715 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 44.8 5.74 ;
      LAYER VIA12 ;
      RECT  43.83 5.47 44.09 5.73 ;
      RECT  44.39 5.47 44.65 5.73 ;
      RECT  41.59 5.47 41.85 5.73 ;
      RECT  38.79 5.47 39.05 5.73 ;
      RECT  37.11 5.47 37.37 5.73 ;
      RECT  34.31 5.47 34.57 5.73 ;
      RECT  32.63 5.47 32.89 5.73 ;
      RECT  28.15 5.47 28.41 5.73 ;
      RECT  28.71 5.47 28.97 5.73 ;
      RECT  29.27 5.47 29.53 5.73 ;
      RECT  29.83 5.47 30.09 5.73 ;
      RECT  25.35 5.47 25.61 5.73 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  44.24 -0.14 44.97 0.14 ;
      RECT  41.325 -0.14 42.73 0.14 ;
      RECT  41.325 0.14 41.555 0.7 ;
      RECT  38.64 -0.14 39.315 0.14 ;
      RECT  39.085 0.14 39.315 0.7 ;
      RECT  36.845 -0.14 37.52 0.14 ;
      RECT  36.845 0.14 37.075 0.7 ;
      RECT  32.365 -0.14 34.835 0.14 ;
      RECT  32.365 0.14 32.595 0.7 ;
      RECT  34.605 0.14 34.835 0.7 ;
      RECT  29.68 -0.14 30.355 0.14 ;
      RECT  30.125 0.14 30.355 0.7 ;
      RECT  25.645 -0.14 28.115 0.14 ;
      RECT  25.645 0.14 25.875 0.7 ;
      RECT  27.885 0.14 28.115 0.7 ;
      RECT  17.36 -0.14 18.48 0.14 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 44.8 0.14 ;
      LAYER VIA12 ;
      RECT  44.39 -0.13 44.65 0.13 ;
      RECT  41.59 -0.13 41.85 0.13 ;
      RECT  42.15 -0.13 42.41 0.13 ;
      RECT  38.79 -0.13 39.05 0.13 ;
      RECT  37.11 -0.13 37.37 0.13 ;
      RECT  32.63 -0.13 32.89 0.13 ;
      RECT  33.19 -0.13 33.45 0.13 ;
      RECT  33.75 -0.13 34.01 0.13 ;
      RECT  34.31 -0.13 34.57 0.13 ;
      RECT  29.83 -0.13 30.09 0.13 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  27.03 -0.13 27.29 0.13 ;
      RECT  27.59 -0.13 27.85 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  18.07 -0.13 18.33 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  24.51 0.98 25.2 1.055 ;
      RECT  24.51 1.055 43.49 1.795 ;
      RECT  42.75 1.795 43.49 3.17 ;
      RECT  42.75 3.17 44.39 3.19 ;
      RECT  42.75 3.19 44.565 3.295 ;
      RECT  9.195 3.295 44.565 3.53 ;
      RECT  9.195 3.53 44.39 3.55 ;
      RECT  9.195 3.55 43.49 4.035 ;
    END
    ANTENNADIFFAREA 38.56 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.98 0.37 7.45 0.6 ;
      RECT  41.82 0.37 44.4 0.6 ;
      RECT  4.66 1.565 9.075 1.795 ;
      RECT  8.845 1.795 9.075 2.405 ;
      RECT  6.605 1.795 6.835 3.805 ;
      RECT  8.845 2.405 42.17 2.635 ;
      RECT  0.18 3.805 8.78 4.035 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
  END
END MDN_BUF_AS_16
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_AS_2
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_AS_2
  CLASS CORE ;
  FOREIGN MDN_BUF_AS_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 1.565 2.06 1.795 ;
      RECT  1.54 1.795 1.82 2.13 ;
      RECT  1.54 2.13 3.81 2.36 ;
      RECT  2.66 2.125 2.94 2.13 ;
      RECT  3.5 2.36 3.81 2.62 ;
      RECT  1.54 2.36 1.82 2.915 ;
      RECT  2.66 2.36 2.94 2.915 ;
    END
    ANTENNADIFFAREA 0.614 ;
    ANTENNAGATEAREA 1.701 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  -0.17 5.46 0.56 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 6.89 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 6.835 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  4.66 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 4.82 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 8.57 0.6 ;
      RECT  3.96 1.565 4.3 1.795 ;
      RECT  4.07 1.795 4.3 2.39 ;
      RECT  4.07 2.39 6.21 2.62 ;
      RECT  4.07 2.62 4.3 3.245 ;
      RECT  2.41 3.245 4.3 3.475 ;
  END
END MDN_BUF_AS_2
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_AS_3
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_AS_3
  CLASS CORE ;
  FOREIGN MDN_BUF_AS_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 1.565 2.06 1.795 ;
      RECT  1.54 1.795 1.82 2.125 ;
      RECT  1.54 2.125 3.81 2.355 ;
      RECT  3.5 2.355 3.81 2.65 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNADIFFAREA 0.614 ;
    ANTENNAGATEAREA 1.701 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  -0.17 5.46 0.56 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 11.37 0.14 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 9.54 1.795 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  4.65 3.245 11.02 3.475 ;
    END
    ANTENNADIFFAREA 7.23 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 9.69 0.6 ;
      RECT  3.96 1.565 4.3 1.795 ;
      RECT  4.07 1.795 4.3 2.39 ;
      RECT  4.07 2.39 8.44 2.62 ;
      RECT  4.07 2.62 4.3 3.245 ;
      RECT  2.38 3.245 4.3 3.475 ;
      RECT  9.35 2.405 10.61 2.635 ;
  END
END MDN_BUF_AS_3
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_AS_4
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_AS_4
  CLASS CORE ;
  FOREIGN MDN_BUF_AS_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 1.565 2.06 1.795 ;
      RECT  1.54 1.795 1.82 2.125 ;
      RECT  1.54 2.125 3.81 2.355 ;
      RECT  3.5 2.355 3.81 2.62 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNADIFFAREA 0.614 ;
    ANTENNAGATEAREA 1.701 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  -0.17 5.46 0.56 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.14 1.565 13.26 1.795 ;
      RECT  11.085 1.795 11.315 3.245 ;
      RECT  4.66 3.245 13.26 3.475 ;
    END
    ANTENNADIFFAREA 9.64 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 11.93 0.6 ;
      RECT  3.96 1.565 4.3 1.795 ;
      RECT  4.07 1.795 4.3 2.39 ;
      RECT  4.07 2.39 10.81 2.62 ;
      RECT  8.235 2.385 8.575 2.39 ;
      RECT  4.07 2.62 4.3 3.245 ;
      RECT  2.38 3.245 4.3 3.475 ;
      RECT  11.59 2.39 13.05 2.62 ;
  END
END MDN_BUF_AS_4
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_AS_6
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_AS_6
  CLASS CORE ;
  FOREIGN MDN_BUF_AS_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.125 ;
      RECT  0.42 2.125 3.81 2.355 ;
      RECT  3.46 2.355 3.81 2.62 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNADIFFAREA 0.614 ;
    ANTENNAGATEAREA 2.268 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.895 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.895 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.705 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.38 1.565 17.74 1.795 ;
      RECT  15.56 1.795 15.79 3.245 ;
      RECT  4.66 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 14.46 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  14.95 0.37 16.41 0.6 ;
      RECT  2.385 1.565 4.325 1.795 ;
      RECT  4.095 1.795 4.325 2.39 ;
      RECT  4.095 2.39 15.29 2.62 ;
      RECT  4.865 2.385 5.205 2.39 ;
      RECT  5.985 2.385 6.325 2.39 ;
      RECT  7.11 2.385 7.45 2.39 ;
      RECT  8.225 2.385 8.565 2.39 ;
      RECT  10.465 2.385 10.805 2.39 ;
      RECT  12.705 2.385 13.045 2.39 ;
      RECT  4.095 2.62 4.325 3.805 ;
      RECT  0.155 3.805 4.325 4.035 ;
      RECT  16.07 2.39 17.53 2.62 ;
  END
END MDN_BUF_AS_6
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_AS_8
#      Description : Non-inverting buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_AS_8
  CLASS CORE ;
  FOREIGN MDN_BUF_AS_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 24.64 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 1.565 2.06 1.795 ;
      RECT  1.54 1.795 1.82 2.125 ;
      RECT  1.54 2.125 6.05 2.355 ;
      RECT  5.79 2.355 6.05 2.62 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
    END
    ANTENNADIFFAREA 0.614 ;
    ANTENNAGATEAREA 2.835 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.81 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  20.72 5.46 21.395 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  -0.17 5.46 0.65 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 24.64 5.74 ;
      LAYER VIA12 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  24.23 5.47 24.49 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 -0.14 24.81 0.14 ;
      RECT  23.405 0.14 23.635 0.67 ;
      RECT  20.72 -0.14 21.395 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  12.205 -0.14 14.675 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 0.65 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 24.64 0.14 ;
      LAYER VIA12 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  20.87 -0.13 21.13 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.86 1.495 24.46 1.865 ;
      RECT  23.405 1.865 23.635 3.175 ;
      RECT  6.9 3.175 24.46 3.545 ;
    END
    ANTENNADIFFAREA 19.28 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  23.91 0.37 24.25 0.6 ;
      RECT  23.91 0.6 24.14 0.9 ;
      RECT  22.79 0.37 23.13 0.6 ;
      RECT  22.9 0.6 23.13 0.9 ;
      RECT  22.9 0.9 24.14 1.13 ;
      RECT  4.66 1.565 6.565 1.795 ;
      RECT  6.335 1.795 6.565 2.405 ;
      RECT  6.335 2.405 23.13 2.635 ;
      RECT  6.335 2.635 6.565 3.805 ;
      RECT  2.42 3.805 6.565 4.035 ;
  END
END MDN_BUF_AS_8
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_S_1
#      Description : Symmetric rise/fall time buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_S_1
  CLASS CORE ;
  FOREIGN MDN_BUF_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.41 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 3.245 ;
      RECT  2.42 3.245 4.3 3.475 ;
    END
    ANTENNADIFFAREA 2.41 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.39 ;
      RECT  1.565 2.39 2.9 2.62 ;
      RECT  1.565 2.62 1.795 3.245 ;
      RECT  0.18 3.245 2.06 3.475 ;
      RECT  0.5 4.365 1.73 4.595 ;
      RECT  0.5 4.595 0.73 5.0 ;
      RECT  1.5 4.595 1.73 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  1.5 5.0 1.85 5.23 ;
      RECT  2.76 4.365 3.945 4.595 ;
      RECT  2.76 4.595 2.99 5.0 ;
      RECT  3.715 4.595 3.945 5.0 ;
      RECT  2.63 5.0 2.99 5.23 ;
      RECT  3.715 5.0 4.09 5.23 ;
  END
END MDN_BUF_S_1
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_S_12
#      Description : Symmetric rise/fall time buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_S_12
  CLASS CORE ;
  FOREIGN MDN_BUF_S_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 33.6 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 6.05 2.355 ;
      RECT  5.74 2.355 6.05 2.62 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  32.365 4.87 32.595 5.46 ;
      RECT  32.365 5.46 33.77 5.74 ;
      RECT  30.125 4.93 30.355 5.46 ;
      RECT  30.125 5.46 30.8 5.74 ;
      RECT  27.885 4.93 28.115 5.46 ;
      RECT  27.44 5.46 28.115 5.74 ;
      RECT  25.645 4.93 25.875 5.46 ;
      RECT  25.2 5.46 25.875 5.74 ;
      RECT  23.405 4.93 23.635 5.46 ;
      RECT  22.96 5.46 23.635 5.74 ;
      RECT  18.925 4.93 19.155 5.46 ;
      RECT  18.925 5.46 21.395 5.74 ;
      RECT  21.165 4.93 21.395 5.46 ;
      RECT  16.685 4.93 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  14.445 4.93 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  9.965 4.93 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.93 12.435 5.46 ;
      RECT  7.725 4.93 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 33.6 5.74 ;
      LAYER VIA12 ;
      RECT  32.63 5.47 32.89 5.73 ;
      RECT  33.19 5.47 33.45 5.73 ;
      RECT  30.39 5.47 30.65 5.73 ;
      RECT  27.59 5.47 27.85 5.73 ;
      RECT  25.35 5.47 25.61 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  20.31 5.47 20.57 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  32.365 -0.14 33.77 0.14 ;
      RECT  32.365 0.14 32.595 0.7 ;
      RECT  30.125 -0.14 30.8 0.14 ;
      RECT  30.125 0.14 30.355 0.7 ;
      RECT  27.44 -0.14 28.115 0.14 ;
      RECT  27.885 0.14 28.115 0.7 ;
      RECT  25.645 -0.14 26.32 0.14 ;
      RECT  25.645 0.14 25.875 0.7 ;
      RECT  23.405 -0.14 24.08 0.14 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  19.99 -0.14 21.395 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  10.64 -0.14 11.37 0.14 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.705 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.695 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 33.6 0.14 ;
      LAYER VIA12 ;
      RECT  32.63 -0.13 32.89 0.13 ;
      RECT  33.19 -0.13 33.45 0.13 ;
      RECT  30.39 -0.13 30.65 0.13 ;
      RECT  27.59 -0.13 27.85 0.13 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  20.31 -0.13 20.57 0.13 ;
      RECT  20.87 -0.13 21.13 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.835 1.515 33.42 1.845 ;
      RECT  19.835 1.845 20.485 3.08 ;
      RECT  26.6 1.845 27.16 3.195 ;
      RECT  6.955 3.08 20.485 3.195 ;
      RECT  6.955 3.195 33.42 3.525 ;
      RECT  6.955 3.525 20.485 3.64 ;
    END
    ANTENNADIFFAREA 28.92 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  19.43 0.37 20.89 0.6 ;
      RECT  26.15 0.37 27.61 0.6 ;
      RECT  3.905 1.565 6.64 1.795 ;
      RECT  6.41 1.795 6.64 2.405 ;
      RECT  6.41 2.405 19.545 2.635 ;
      RECT  6.41 2.635 6.64 3.245 ;
      RECT  6.045 3.245 6.64 3.475 ;
      RECT  6.045 3.475 6.275 4.365 ;
      RECT  0.17 4.365 6.275 4.595 ;
      RECT  20.775 2.405 26.265 2.635 ;
      RECT  27.495 2.405 33.21 2.635 ;
  END
END MDN_BUF_S_12
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_S_16
#      Description : Symmetric rise/fall time buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_S_16
  CLASS CORE ;
  FOREIGN MDN_BUF_S_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 44.8 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 8.31 2.355 ;
      RECT  8.03 2.355 8.31 2.695 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
    END
    ANTENNAGATEAREA 4.536 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  43.565 4.87 43.795 5.46 ;
      RECT  43.565 5.46 44.97 5.74 ;
      RECT  41.325 4.93 41.555 5.46 ;
      RECT  41.325 5.46 42.56 5.74 ;
      RECT  39.085 4.93 39.315 5.46 ;
      RECT  38.64 5.46 39.315 5.74 ;
      RECT  36.845 4.93 37.075 5.46 ;
      RECT  36.4 5.46 37.075 5.74 ;
      RECT  32.365 4.93 32.595 5.46 ;
      RECT  32.365 5.46 34.835 5.74 ;
      RECT  34.605 4.93 34.835 5.46 ;
      RECT  30.125 4.93 30.355 5.46 ;
      RECT  29.68 5.46 30.355 5.74 ;
      RECT  27.885 4.93 28.115 5.46 ;
      RECT  27.44 5.46 28.115 5.74 ;
      RECT  25.645 4.93 25.875 5.46 ;
      RECT  25.2 5.46 25.875 5.74 ;
      RECT  21.165 4.93 21.395 5.46 ;
      RECT  21.165 5.46 23.635 5.74 ;
      RECT  23.405 4.93 23.635 5.46 ;
      RECT  18.925 4.93 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  16.685 4.93 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  12.205 4.93 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 4.93 14.675 5.46 ;
      RECT  9.965 4.93 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.905 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 44.8 5.74 ;
      LAYER VIA12 ;
      RECT  43.83 5.47 44.09 5.73 ;
      RECT  44.39 5.47 44.65 5.73 ;
      RECT  41.59 5.47 41.85 5.73 ;
      RECT  42.15 5.47 42.41 5.73 ;
      RECT  38.79 5.47 39.05 5.73 ;
      RECT  36.55 5.47 36.81 5.73 ;
      RECT  32.63 5.47 32.89 5.73 ;
      RECT  33.19 5.47 33.45 5.73 ;
      RECT  33.75 5.47 34.01 5.73 ;
      RECT  34.31 5.47 34.57 5.73 ;
      RECT  29.83 5.47 30.09 5.73 ;
      RECT  27.59 5.47 27.85 5.73 ;
      RECT  25.35 5.47 25.61 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  22.55 5.47 22.81 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  43.565 -0.14 44.97 0.14 ;
      RECT  43.565 0.14 43.795 0.7 ;
      RECT  41.325 -0.14 42.0 0.14 ;
      RECT  41.325 0.14 41.555 0.7 ;
      RECT  38.64 -0.14 39.315 0.14 ;
      RECT  39.085 0.14 39.315 0.7 ;
      RECT  36.4 -0.14 37.075 0.14 ;
      RECT  36.845 0.14 37.075 0.7 ;
      RECT  32.365 -0.14 34.835 0.14 ;
      RECT  32.365 0.14 32.595 0.7 ;
      RECT  34.605 0.14 34.835 0.7 ;
      RECT  29.68 -0.14 30.355 0.14 ;
      RECT  30.125 0.14 30.355 0.7 ;
      RECT  27.44 -0.14 28.115 0.14 ;
      RECT  27.885 0.14 28.115 0.7 ;
      RECT  21.84 -0.14 22.57 0.14 ;
      RECT  12.88 -0.14 13.61 0.14 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.705 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 44.8 0.14 ;
      LAYER VIA12 ;
      RECT  43.83 -0.13 44.09 0.13 ;
      RECT  44.39 -0.13 44.65 0.13 ;
      RECT  41.59 -0.13 41.85 0.13 ;
      RECT  38.79 -0.13 39.05 0.13 ;
      RECT  36.55 -0.13 36.81 0.13 ;
      RECT  32.63 -0.13 32.89 0.13 ;
      RECT  33.19 -0.13 33.45 0.13 ;
      RECT  33.75 -0.13 34.01 0.13 ;
      RECT  34.31 -0.13 34.57 0.13 ;
      RECT  29.83 -0.13 30.09 0.13 ;
      RECT  27.59 -0.13 27.85 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  26.81 1.005 43.205 1.01 ;
      RECT  26.465 1.01 43.205 1.125 ;
      RECT  26.465 1.125 43.21 1.565 ;
      RECT  26.465 1.565 44.62 1.745 ;
      RECT  42.18 1.745 44.62 1.795 ;
      RECT  26.465 1.745 27.295 3.045 ;
      RECT  42.18 1.795 43.21 1.82 ;
      RECT  42.37 1.82 43.21 3.045 ;
      RECT  9.195 3.045 43.21 3.245 ;
      RECT  9.195 3.245 44.62 3.475 ;
      RECT  9.195 3.475 43.21 3.55 ;
      RECT  9.195 3.55 43.205 3.785 ;
    END
    ANTENNADIFFAREA 38.56 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  26.15 0.37 27.61 0.6 ;
      RECT  4.66 1.565 8.91 1.795 ;
      RECT  8.68 1.795 8.91 2.39 ;
      RECT  8.68 2.39 26.21 2.62 ;
      RECT  25.98 2.335 26.21 2.39 ;
      RECT  25.98 2.62 26.21 2.675 ;
      RECT  8.68 2.62 8.91 3.245 ;
      RECT  8.285 3.245 8.91 3.475 ;
      RECT  8.285 3.475 8.515 3.805 ;
      RECT  0.18 3.805 8.515 4.035 ;
      RECT  27.55 2.335 27.78 2.39 ;
      RECT  27.55 2.39 41.945 2.62 ;
      RECT  27.55 2.62 27.78 2.675 ;
      RECT  43.08 4.365 44.255 4.595 ;
      RECT  43.08 4.595 43.31 5.0 ;
      RECT  44.025 4.595 44.255 5.0 ;
      RECT  41.83 5.0 43.31 5.23 ;
      RECT  44.025 5.0 44.41 5.23 ;
  END
END MDN_BUF_S_16
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_S_2
#      Description : Symmetric rise/fall time buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_S_2
  CLASS CORE ;
  FOREIGN MDN_BUF_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.41 1.565 5.715 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  2.42 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 4.82 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.775 1.575 2.005 2.39 ;
      RECT  1.775 2.39 5.21 2.62 ;
      RECT  1.775 2.62 2.005 3.245 ;
      RECT  0.18 3.245 2.005 3.475 ;
      RECT  0.52 4.365 1.695 4.595 ;
      RECT  0.52 4.595 0.75 5.0 ;
      RECT  1.465 4.595 1.695 5.0 ;
      RECT  0.39 5.0 0.75 5.23 ;
      RECT  1.465 5.0 1.85 5.23 ;
      RECT  5.0 4.365 6.2 4.595 ;
      RECT  5.0 4.595 5.23 5.0 ;
      RECT  5.97 4.595 6.2 5.0 ;
      RECT  4.87 5.0 5.23 5.23 ;
      RECT  5.97 5.0 6.315 5.23 ;
  END
END MDN_BUF_S_2
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_S_3
#      Description : Symmetric rise/fall time buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_S_3
  CLASS CORE ;
  FOREIGN MDN_BUF_S_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.17 1.565 8.78 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  2.42 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 7.23 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.39 ;
      RECT  1.565 2.39 7.395 2.62 ;
      RECT  1.565 2.62 1.795 3.245 ;
      RECT  0.18 3.245 2.06 3.475 ;
      RECT  0.52 4.365 1.715 4.595 ;
      RECT  0.52 4.595 0.75 5.0 ;
      RECT  1.485 4.595 1.715 5.0 ;
      RECT  0.39 5.0 0.75 5.23 ;
      RECT  1.485 5.0 1.85 5.23 ;
      RECT  7.24 4.365 8.425 4.595 ;
      RECT  7.24 4.595 7.47 5.0 ;
      RECT  8.195 4.595 8.425 5.0 ;
      RECT  7.11 5.0 7.47 5.23 ;
      RECT  8.195 5.0 8.57 5.23 ;
  END
END MDN_BUF_S_3
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_S_4
#      Description : Symmetric rise/fall time buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_S_4
  CLASS CORE ;
  FOREIGN MDN_BUF_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.555 1.565 11.02 1.795 ;
      RECT  6.555 1.795 7.09 1.82 ;
      RECT  6.555 1.82 6.885 3.22 ;
      RECT  6.35 3.22 7.09 3.245 ;
      RECT  2.42 3.245 11.02 3.475 ;
    END
    ANTENNADIFFAREA 9.64 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.39 ;
      RECT  1.565 2.39 6.305 2.62 ;
      RECT  1.565 2.62 1.795 3.245 ;
      RECT  0.18 3.245 2.06 3.475 ;
      RECT  7.13 2.39 10.81 2.62 ;
      RECT  0.52 4.365 1.695 4.595 ;
      RECT  0.52 4.595 0.75 5.0 ;
      RECT  1.465 4.595 1.695 5.0 ;
      RECT  0.39 5.0 0.75 5.23 ;
      RECT  1.465 5.0 1.85 5.23 ;
  END
END MDN_BUF_S_4
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_S_6
#      Description : Symmetric rise/fall time buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_S_6
  CLASS CORE ;
  FOREIGN MDN_BUF_S_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.035 2.355 ;
      RECT  3.805 2.355 4.035 2.67 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 18.09 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  11.76 -0.14 12.435 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  8.79 -0.14 9.52 0.14 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.035 1.54 17.735 1.565 ;
      RECT  11.035 1.565 17.74 1.795 ;
      RECT  11.035 1.795 17.735 1.87 ;
      RECT  11.035 1.87 11.365 3.73 ;
      RECT  10.825 3.73 17.74 3.805 ;
      RECT  4.66 3.805 17.74 4.035 ;
      RECT  10.825 4.035 17.74 4.06 ;
    END
    ANTENNADIFFAREA 14.46 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 11.93 0.6 ;
      RECT  2.42 1.565 4.595 1.795 ;
      RECT  4.365 1.795 4.595 2.39 ;
      RECT  4.365 2.39 10.66 2.62 ;
      RECT  5.995 2.385 6.335 2.39 ;
      RECT  7.11 2.385 7.45 2.39 ;
      RECT  8.23 2.385 8.57 2.39 ;
      RECT  9.35 2.385 9.69 2.39 ;
      RECT  4.365 2.62 4.595 3.07 ;
      RECT  3.805 3.07 4.595 3.3 ;
      RECT  3.805 3.3 4.035 3.805 ;
      RECT  0.18 3.805 4.035 4.035 ;
      RECT  11.76 2.39 17.42 2.62 ;
      RECT  14.94 5.0 16.41 5.23 ;
  END
END MDN_BUF_S_6
#-----------------------------------------------------------------------
#      Cell        : MDN_BUF_S_8
#      Description : Symmetric rise/fall time buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUF_S_8
  CLASS CORE ;
  FOREIGN MDN_BUF_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 3.81 2.355 ;
      RECT  3.55 2.355 3.81 2.69 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 22.57 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  7.725 4.895 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  20.31 5.47 20.57 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.925 -0.14 19.6 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  13.27 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.205 1.49 22.165 1.96 ;
      RECT  13.205 1.96 13.675 3.08 ;
      RECT  4.715 3.08 22.155 3.19 ;
      RECT  4.715 3.19 22.165 3.53 ;
      RECT  4.715 3.53 22.155 3.55 ;
    END
    ANTENNADIFFAREA 19.28 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  21.67 0.37 22.01 0.6 ;
      RECT  21.67 0.6 21.9 1.005 ;
      RECT  20.55 0.37 20.89 0.6 ;
      RECT  20.66 0.6 20.89 1.005 ;
      RECT  19.43 0.37 19.77 0.6 ;
      RECT  19.43 0.6 19.66 1.005 ;
      RECT  18.31 0.37 18.65 0.6 ;
      RECT  18.42 0.6 18.65 1.005 ;
      RECT  17.19 0.37 17.53 0.6 ;
      RECT  17.19 0.6 17.42 1.005 ;
      RECT  16.07 0.37 16.41 0.6 ;
      RECT  16.18 0.6 16.41 1.005 ;
      RECT  14.95 0.37 15.29 0.6 ;
      RECT  14.95 0.6 15.18 1.005 ;
      RECT  12.68 0.37 14.17 0.6 ;
      RECT  13.94 0.6 14.17 1.005 ;
      RECT  12.68 0.6 12.91 2.405 ;
      RECT  13.94 1.005 21.9 1.235 ;
      RECT  2.42 1.565 4.3 1.795 ;
      RECT  4.07 1.795 4.3 2.405 ;
      RECT  4.07 2.405 12.91 2.635 ;
      RECT  4.07 2.635 4.3 3.035 ;
      RECT  3.805 3.035 4.3 3.265 ;
      RECT  3.805 3.265 4.035 3.805 ;
      RECT  0.175 3.805 4.035 4.035 ;
  END
END MDN_BUF_S_8
#-----------------------------------------------------------------------
#      Cell        : MDN_BUFTS_1
#      Description : Internal tri-state buffer (active hi-enable)
#      Equation    : X=tristate(enable=EN,data=A)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUFTS_1
  CLASS CORE ;
  FOREIGN MDN_BUFTS_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 4.365 6.275 4.595 ;
      RECT  3.805 4.595 4.035 5.0 ;
      RECT  6.045 4.595 6.275 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
      RECT  5.99 5.0 6.33 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.925 0.6 5.155 1.005 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  1.565 1.005 5.155 1.235 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  2.42 4.365 2.915 4.595 ;
      RECT  2.685 4.595 2.915 5.46 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  1.005 5.46 2.915 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 0.14 5.715 1.565 ;
      RECT  4.66 1.565 5.715 1.795 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 7.955 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  7.725 3.245 8.785 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 8.57 0.6 ;
      RECT  8.245 0.6 8.475 1.005 ;
      RECT  6.045 1.005 8.475 1.235 ;
      RECT  6.045 1.235 6.275 1.565 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 3.245 ;
      RECT  4.66 3.245 6.54 3.475 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.39 ;
      RECT  1.565 2.39 2.765 2.62 ;
      RECT  1.565 2.62 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  2.42 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 3.805 ;
      RECT  3.805 3.805 7.395 4.035 ;
      RECT  7.165 2.33 7.395 3.805 ;
  END
END MDN_BUFTS_1
#-----------------------------------------------------------------------
#      Cell        : MDN_BUFTS_12
#      Description : Internal tri-state buffer (active hi-enable)
#      Equation    : X=tristate(enable=EN,data=A)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUFTS_12
  CLASS CORE ;
  FOREIGN MDN_BUFTS_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 44.8 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 16.38 2.355 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 3.85 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.5 2.355 3.85 2.94 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  43.565 4.9 43.795 5.46 ;
      RECT  43.565 5.46 44.97 5.74 ;
      RECT  39.085 4.9 39.315 5.46 ;
      RECT  39.085 5.46 41.555 5.74 ;
      RECT  41.325 4.9 41.555 5.46 ;
      RECT  34.605 4.9 34.835 5.46 ;
      RECT  34.605 5.46 37.075 5.74 ;
      RECT  36.845 4.9 37.075 5.46 ;
      RECT  30.125 4.9 30.355 5.46 ;
      RECT  30.125 5.46 32.595 5.74 ;
      RECT  32.365 4.9 32.595 5.46 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.645 5.46 28.115 5.74 ;
      RECT  27.885 4.9 28.115 5.46 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 23.635 5.74 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  14.445 4.87 14.675 5.46 ;
      RECT  14.445 5.46 16.915 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 5.715 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 44.8 5.74 ;
      LAYER VIA12 ;
      RECT  43.83 5.47 44.09 5.73 ;
      RECT  44.39 5.47 44.65 5.73 ;
      RECT  39.35 5.47 39.61 5.73 ;
      RECT  39.91 5.47 40.17 5.73 ;
      RECT  40.47 5.47 40.73 5.73 ;
      RECT  41.03 5.47 41.29 5.73 ;
      RECT  34.87 5.47 35.13 5.73 ;
      RECT  35.43 5.47 35.69 5.73 ;
      RECT  35.99 5.47 36.25 5.73 ;
      RECT  36.55 5.47 36.81 5.73 ;
      RECT  30.39 5.47 30.65 5.73 ;
      RECT  30.95 5.47 31.21 5.73 ;
      RECT  31.51 5.47 31.77 5.73 ;
      RECT  32.07 5.47 32.33 5.73 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  27.03 5.47 27.29 5.73 ;
      RECT  27.59 5.47 27.85 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  22.55 5.47 22.81 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  43.565 -0.14 44.97 0.14 ;
      RECT  43.565 0.14 43.795 0.73 ;
      RECT  39.085 -0.14 41.555 0.14 ;
      RECT  39.085 0.14 39.315 0.73 ;
      RECT  41.325 0.14 41.555 0.73 ;
      RECT  34.605 -0.14 37.075 0.14 ;
      RECT  34.605 0.14 34.835 0.73 ;
      RECT  36.845 0.14 37.075 0.73 ;
      RECT  30.125 -0.14 32.595 0.14 ;
      RECT  32.365 0.14 32.595 0.675 ;
      RECT  30.125 0.14 30.355 0.73 ;
      RECT  25.645 -0.14 28.115 0.14 ;
      RECT  25.645 0.14 25.875 0.73 ;
      RECT  27.885 0.14 28.115 0.73 ;
      RECT  21.165 -0.14 23.635 0.14 ;
      RECT  21.165 0.14 21.395 0.73 ;
      RECT  23.405 0.14 23.635 0.73 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  11.76 -0.14 12.435 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  7.725 -0.14 10.195 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 44.8 0.14 ;
      LAYER VIA12 ;
      RECT  43.83 -0.13 44.09 0.13 ;
      RECT  44.39 -0.13 44.65 0.13 ;
      RECT  39.35 -0.13 39.61 0.13 ;
      RECT  39.91 -0.13 40.17 0.13 ;
      RECT  40.47 -0.13 40.73 0.13 ;
      RECT  41.03 -0.13 41.29 0.13 ;
      RECT  34.87 -0.13 35.13 0.13 ;
      RECT  35.43 -0.13 35.69 0.13 ;
      RECT  35.99 -0.13 36.25 0.13 ;
      RECT  36.55 -0.13 36.81 0.13 ;
      RECT  30.39 -0.13 30.65 0.13 ;
      RECT  30.95 -0.13 31.21 0.13 ;
      RECT  31.51 -0.13 31.77 0.13 ;
      RECT  32.07 -0.13 32.33 0.13 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  27.03 -0.13 27.29 0.13 ;
      RECT  27.59 -0.13 27.85 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  22.55 -0.13 22.81 0.13 ;
      RECT  23.11 -0.13 23.37 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER METAL1 ;
      RECT  18.07 1.465 44.565 2.025 ;
      RECT  44.005 2.025 44.565 2.99 ;
      RECT  19.64 2.99 44.565 3.55 ;
    END
    ANTENNADIFFAREA 18.144 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  44.07 0.37 44.41 0.6 ;
      RECT  44.07 0.6 44.3 1.005 ;
      RECT  41.83 0.37 42.17 0.6 ;
      RECT  41.83 0.6 42.06 1.005 ;
      RECT  39.59 0.37 39.93 0.6 ;
      RECT  39.59 0.6 39.82 1.005 ;
      RECT  37.35 0.37 37.69 0.6 ;
      RECT  37.35 0.6 37.58 1.005 ;
      RECT  35.11 0.37 35.45 0.6 ;
      RECT  35.11 0.6 35.34 1.005 ;
      RECT  32.87 0.37 33.21 0.6 ;
      RECT  32.87 0.6 33.1 1.005 ;
      RECT  30.63 0.37 30.97 0.6 ;
      RECT  30.63 0.6 30.86 1.005 ;
      RECT  28.39 0.37 28.73 0.6 ;
      RECT  28.39 0.6 28.62 1.005 ;
      RECT  26.15 0.37 26.49 0.6 ;
      RECT  26.15 0.6 26.38 1.005 ;
      RECT  23.91 0.37 24.25 0.6 ;
      RECT  23.91 0.6 24.14 1.005 ;
      RECT  21.67 0.37 22.01 0.6 ;
      RECT  21.67 0.6 21.9 1.005 ;
      RECT  19.43 0.37 19.77 0.6 ;
      RECT  19.43 0.6 19.66 1.005 ;
      RECT  13.62 1.005 44.3 1.235 ;
      RECT  16.685 1.235 16.915 3.245 ;
      RECT  15.16 3.245 16.915 3.475 ;
      RECT  12.765 0.445 16.97 0.675 ;
      RECT  12.765 0.675 12.995 1.005 ;
      RECT  0.18 1.005 12.995 1.235 ;
      RECT  3.96 1.565 4.37 1.795 ;
      RECT  4.14 1.795 4.37 2.125 ;
      RECT  4.14 2.125 4.595 2.355 ;
      RECT  4.365 2.355 4.595 2.405 ;
      RECT  4.365 2.405 7.45 2.635 ;
      RECT  4.365 2.635 4.595 3.245 ;
      RECT  3.96 3.245 4.595 3.475 ;
      RECT  17.245 2.405 43.29 2.635 ;
      RECT  17.245 2.635 17.475 3.805 ;
      RECT  4.66 1.565 13.26 1.795 ;
      RECT  9.965 1.795 10.195 3.805 ;
      RECT  9.965 3.805 17.475 4.035 ;
      RECT  4.66 3.805 9.075 4.035 ;
      RECT  8.845 4.035 9.075 4.365 ;
      RECT  8.845 4.365 13.26 4.595 ;
      RECT  13.62 4.365 16.225 4.595 ;
      RECT  13.62 4.595 13.85 4.925 ;
      RECT  0.165 4.365 8.515 4.595 ;
      RECT  8.285 4.595 8.515 4.925 ;
      RECT  8.285 4.925 13.85 5.155 ;
  END
END MDN_BUFTS_12
#-----------------------------------------------------------------------
#      Cell        : MDN_BUFTS_2
#      Description : Internal tri-state buffer (active hi-enable)
#      Equation    : X=tristate(enable=EN,data=A)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUFTS_2
  CLASS CORE ;
  FOREIGN MDN_BUFTS_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 4.365 6.275 4.595 ;
      RECT  3.805 4.595 4.035 5.0 ;
      RECT  6.045 4.595 6.275 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
      RECT  5.99 5.0 6.33 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 0.37 5.21 0.6 ;
      RECT  3.805 0.6 4.035 1.005 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  1.565 1.005 4.035 1.235 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  2.42 4.365 2.915 4.595 ;
      RECT  2.685 4.595 2.915 5.46 ;
      RECT  2.07 5.46 2.915 5.74 ;
      RECT  1.005 4.865 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.485 0.14 5.715 1.005 ;
      RECT  4.66 1.005 5.715 1.235 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.69 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER METAL1 ;
      RECT  6.87 1.565 10.195 1.795 ;
      RECT  9.965 1.795 10.195 3.245 ;
      RECT  8.44 3.245 11.02 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  10.445 0.37 10.81 0.6 ;
      RECT  10.445 0.6 10.675 0.995 ;
      RECT  8.205 0.37 8.57 0.6 ;
      RECT  8.205 0.6 8.435 0.995 ;
      RECT  6.34 0.995 10.675 1.225 ;
      RECT  6.34 1.225 6.57 1.565 ;
      RECT  5.48 1.565 6.57 1.795 ;
      RECT  5.48 1.795 5.71 3.245 ;
      RECT  4.66 3.245 6.555 3.475 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.41 ;
      RECT  1.565 2.41 2.805 2.64 ;
      RECT  1.565 2.64 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  7.16 2.385 9.47 2.615 ;
      RECT  7.16 2.615 7.39 3.805 ;
      RECT  2.39 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 3.805 ;
      RECT  3.805 3.805 7.39 4.035 ;
  END
END MDN_BUFTS_2
#-----------------------------------------------------------------------
#      Cell        : MDN_BUFTS_3
#      Description : Internal tri-state buffer (active hi-enable)
#      Equation    : X=tristate(enable=EN,data=A)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUFTS_3
  CLASS CORE ;
  FOREIGN MDN_BUFTS_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 4.365 6.275 4.595 ;
      RECT  3.805 4.595 4.035 5.0 ;
      RECT  6.045 4.595 6.275 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
      RECT  5.99 5.0 6.33 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 0.37 5.215 0.6 ;
      RECT  3.805 0.6 4.035 1.005 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  1.565 1.005 4.035 1.235 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  2.42 4.365 2.915 4.595 ;
      RECT  2.685 4.595 2.915 5.46 ;
      RECT  2.07 5.46 2.915 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.485 0.14 5.715 1.005 ;
      RECT  4.63 1.005 5.715 1.235 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 12.435 1.795 ;
      RECT  12.205 1.795 12.435 3.245 ;
      RECT  8.44 3.245 13.26 3.475 ;
    END
    ANTENNADIFFAREA 4.536 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  12.665 0.37 13.05 0.6 ;
      RECT  12.665 0.6 12.895 1.005 ;
      RECT  10.47 0.37 10.81 0.6 ;
      RECT  10.47 0.6 10.7 1.005 ;
      RECT  8.23 0.37 8.57 0.6 ;
      RECT  8.23 0.6 8.46 1.005 ;
      RECT  6.31 1.005 12.895 1.235 ;
      RECT  6.31 1.235 6.54 1.565 ;
      RECT  5.485 1.565 6.54 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  4.66 3.245 6.54 3.475 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.42 ;
      RECT  1.565 2.42 2.97 2.65 ;
      RECT  1.565 2.65 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  7.165 2.39 11.885 2.62 ;
      RECT  7.165 2.62 7.395 3.805 ;
      RECT  2.42 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 3.805 ;
      RECT  3.805 3.805 7.395 4.035 ;
  END
END MDN_BUFTS_3
#-----------------------------------------------------------------------
#      Cell        : MDN_BUFTS_4
#      Description : Internal tri-state buffer (active hi-enable)
#      Equation    : X=tristate(enable=EN,data=A)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUFTS_4
  CLASS CORE ;
  FOREIGN MDN_BUFTS_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 4.365 6.275 4.595 ;
      RECT  3.805 4.595 4.035 5.0 ;
      RECT  6.045 4.595 6.275 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
      RECT  5.99 5.0 6.33 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 0.37 5.21 0.6 ;
      RECT  3.805 0.6 4.035 1.005 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  1.565 1.005 4.035 1.235 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  2.42 4.365 2.915 4.595 ;
      RECT  2.685 4.595 2.915 5.46 ;
      RECT  2.07 5.46 2.915 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  5.46 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.46 0.14 5.69 1.005 ;
      RECT  4.63 1.005 5.69 1.235 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 14.675 1.795 ;
      RECT  14.445 1.795 14.675 3.245 ;
      RECT  8.44 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  14.91 0.37 15.29 0.6 ;
      RECT  14.91 0.6 15.14 1.01 ;
      RECT  12.675 0.37 13.05 0.6 ;
      RECT  12.675 0.6 12.905 1.01 ;
      RECT  10.435 0.37 10.81 0.6 ;
      RECT  10.435 0.6 10.665 1.01 ;
      RECT  8.195 0.37 8.57 0.6 ;
      RECT  8.195 0.6 8.425 1.01 ;
      RECT  6.315 1.01 15.14 1.24 ;
      RECT  6.315 1.24 6.545 1.565 ;
      RECT  5.485 1.565 6.545 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  4.655 3.245 6.545 3.475 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.39 ;
      RECT  1.565 2.39 2.78 2.62 ;
      RECT  1.565 2.62 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  7.165 2.405 14.17 2.635 ;
      RECT  7.165 2.635 7.395 3.805 ;
      RECT  2.42 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 3.805 ;
      RECT  3.805 3.805 7.395 4.035 ;
  END
END MDN_BUFTS_4
#-----------------------------------------------------------------------
#      Cell        : MDN_BUFTS_6
#      Description : Internal tri-state buffer (active hi-enable)
#      Equation    : X=tristate(enable=EN,data=A)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUFTS_6
  CLASS CORE ;
  FOREIGN MDN_BUFTS_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 24.64 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 10.605 2.355 ;
      RECT  10.22 2.355 10.605 2.43 ;
      RECT  9.405 2.355 9.635 2.69 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  10.375 2.43 10.605 2.675 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 3.815 2.355 ;
      RECT  3.22 2.355 3.815 2.67 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  3.22 2.67 3.5 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 4.93 23.635 5.46 ;
      RECT  23.405 5.46 24.81 5.74 ;
      RECT  21.165 4.93 21.395 5.46 ;
      RECT  21.165 5.46 21.84 5.74 ;
      RECT  18.925 4.93 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  16.685 4.93 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  12.205 4.93 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 4.93 14.675 5.46 ;
      RECT  9.965 4.935 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  5.485 4.935 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 24.64 5.74 ;
      LAYER VIA12 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  24.23 5.47 24.49 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 -0.14 24.81 0.14 ;
      RECT  23.405 0.14 23.635 0.73 ;
      RECT  21.165 -0.14 21.84 0.14 ;
      RECT  21.165 0.14 21.395 0.73 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  12.205 -0.14 14.675 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 24.64 0.14 ;
      LAYER VIA12 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER METAL1 ;
      RECT  11.38 1.515 23.685 1.845 ;
      RECT  23.355 1.845 23.685 3.195 ;
      RECT  12.92 3.195 24.455 3.245 ;
      RECT  12.92 3.245 24.46 3.475 ;
      RECT  12.92 3.475 24.455 3.525 ;
    END
    ANTENNADIFFAREA 9.072 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  23.865 0.37 24.25 0.6 ;
      RECT  23.865 0.6 24.095 0.97 ;
      RECT  21.625 0.37 22.01 0.6 ;
      RECT  21.625 0.6 21.855 0.97 ;
      RECT  19.385 0.37 19.77 0.6 ;
      RECT  19.385 0.6 19.615 0.97 ;
      RECT  17.145 0.37 17.53 0.6 ;
      RECT  17.145 0.6 17.375 0.97 ;
      RECT  14.905 0.37 15.29 0.6 ;
      RECT  14.905 0.6 15.135 0.97 ;
      RECT  12.665 0.37 13.05 0.6 ;
      RECT  12.665 0.6 12.905 0.97 ;
      RECT  12.665 0.97 24.095 1.005 ;
      RECT  10.85 1.005 24.095 1.235 ;
      RECT  10.85 1.235 11.08 1.565 ;
      RECT  9.14 1.565 11.08 1.795 ;
      RECT  10.85 1.795 11.08 3.03 ;
      RECT  9.11 3.03 11.08 3.26 ;
      RECT  0.18 1.005 10.25 1.235 ;
      RECT  3.96 1.565 4.36 1.795 ;
      RECT  4.13 1.795 4.36 2.39 ;
      RECT  4.13 2.39 6.125 2.62 ;
      RECT  4.365 2.62 4.595 3.245 ;
      RECT  3.915 3.245 4.595 3.475 ;
      RECT  11.645 2.405 22.94 2.635 ;
      RECT  11.645 2.635 11.875 3.805 ;
      RECT  4.66 1.565 8.8 1.795 ;
      RECT  6.605 1.795 6.835 3.555 ;
      RECT  6.605 3.555 9.635 3.785 ;
      RECT  9.405 3.785 9.635 3.805 ;
      RECT  9.405 3.805 11.875 4.035 ;
      RECT  4.66 4.015 8.78 4.245 ;
      RECT  0.15 4.365 4.36 4.475 ;
      RECT  0.15 4.475 11.02 4.595 ;
      RECT  4.13 4.595 11.02 4.705 ;
      RECT  10.68 4.705 11.02 4.71 ;
  END
END MDN_BUFTS_6
#-----------------------------------------------------------------------
#      Cell        : MDN_BUFTS_8
#      Description : Internal tri-state buffer (active hi-enable)
#      Equation    : X=tristate(enable=EN,data=A)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUFTS_8
  CLASS CORE ;
  FOREIGN MDN_BUFTS_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 29.12 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 10.78 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 4.06 2.355 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  27.885 4.9 28.115 5.46 ;
      RECT  27.885 5.46 29.29 5.74 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.2 5.46 25.875 5.74 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  22.96 5.46 23.635 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 21.84 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  0.445 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 29.12 5.74 ;
      LAYER VIA12 ;
      RECT  28.15 5.47 28.41 5.73 ;
      RECT  28.71 5.47 28.97 5.73 ;
      RECT  25.35 5.47 25.61 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  27.885 -0.14 29.29 0.14 ;
      RECT  27.885 0.14 28.115 0.7 ;
      RECT  25.2 -0.14 25.875 0.14 ;
      RECT  25.645 0.14 25.875 0.7 ;
      RECT  23.405 -0.14 24.08 0.14 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  21.165 -0.14 21.84 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  12.205 -0.14 14.675 0.14 ;
      RECT  12.205 0.14 12.435 0.52 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.445 1.005 2.06 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 29.12 0.14 ;
      LAYER VIA12 ;
      RECT  28.15 -0.13 28.41 0.13 ;
      RECT  28.71 -0.13 28.97 0.13 ;
      RECT  25.35 -0.13 25.61 0.13 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER METAL1 ;
      RECT  11.16 1.205 11.665 1.21 ;
      RECT  11.16 1.21 11.875 1.435 ;
      RECT  11.38 1.435 11.875 1.44 ;
      RECT  11.57 1.44 11.875 1.495 ;
      RECT  11.57 1.495 28.745 1.54 ;
      RECT  11.645 1.54 28.745 1.865 ;
      RECT  28.375 1.865 28.745 3.175 ;
      RECT  12.975 3.175 28.885 3.545 ;
    END
    ANTENNADIFFAREA 12.096 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  28.39 0.37 28.945 0.6 ;
      RECT  28.715 0.6 28.945 1.005 ;
      RECT  26.15 0.37 26.49 0.6 ;
      RECT  26.15 0.6 26.38 1.005 ;
      RECT  23.91 0.37 24.25 0.6 ;
      RECT  23.91 0.6 24.14 1.005 ;
      RECT  21.67 0.37 22.01 0.6 ;
      RECT  21.67 0.6 21.9 1.005 ;
      RECT  19.43 0.37 19.77 0.6 ;
      RECT  19.43 0.6 19.66 1.005 ;
      RECT  17.19 0.37 17.53 0.6 ;
      RECT  17.19 0.6 17.42 1.005 ;
      RECT  14.95 0.37 15.29 0.6 ;
      RECT  14.95 0.6 15.18 1.005 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 0.75 ;
      RECT  10.525 0.445 11.77 0.45 ;
      RECT  10.525 0.45 11.775 0.455 ;
      RECT  10.525 0.455 11.78 0.46 ;
      RECT  10.525 0.46 11.785 0.465 ;
      RECT  10.525 0.465 11.79 0.47 ;
      RECT  10.525 0.47 11.795 0.475 ;
      RECT  10.525 0.475 11.8 0.48 ;
      RECT  10.525 0.48 11.805 0.485 ;
      RECT  10.525 0.485 11.81 0.49 ;
      RECT  10.525 0.49 11.815 0.495 ;
      RECT  10.525 0.495 11.82 0.5 ;
      RECT  10.525 0.5 11.825 0.505 ;
      RECT  10.525 0.505 11.83 0.51 ;
      RECT  10.525 0.51 11.835 0.515 ;
      RECT  10.525 0.515 11.84 0.52 ;
      RECT  10.525 0.52 11.845 0.525 ;
      RECT  10.525 0.525 11.85 0.53 ;
      RECT  10.525 0.53 11.855 0.535 ;
      RECT  10.525 0.535 11.86 0.54 ;
      RECT  10.525 0.54 11.865 0.545 ;
      RECT  10.525 0.545 11.87 0.55 ;
      RECT  10.525 0.55 11.875 0.555 ;
      RECT  10.525 0.555 11.88 0.56 ;
      RECT  10.525 0.56 11.885 0.565 ;
      RECT  10.525 0.565 11.89 0.57 ;
      RECT  10.525 0.57 11.895 0.575 ;
      RECT  10.525 0.575 11.9 0.58 ;
      RECT  10.525 0.58 11.905 0.585 ;
      RECT  10.525 0.585 11.91 0.59 ;
      RECT  10.525 0.59 11.915 0.595 ;
      RECT  10.525 0.595 11.92 0.6 ;
      RECT  10.525 0.6 11.925 0.605 ;
      RECT  10.525 0.605 11.93 0.61 ;
      RECT  10.525 0.61 11.935 0.615 ;
      RECT  10.525 0.615 11.94 0.62 ;
      RECT  10.525 0.62 11.945 0.625 ;
      RECT  10.525 0.625 11.95 0.63 ;
      RECT  10.525 0.63 11.955 0.635 ;
      RECT  10.525 0.635 11.96 0.64 ;
      RECT  10.525 0.64 11.965 0.645 ;
      RECT  10.525 0.645 11.97 0.65 ;
      RECT  10.525 0.65 11.975 0.655 ;
      RECT  10.525 0.655 11.98 0.66 ;
      RECT  10.525 0.66 11.985 0.665 ;
      RECT  10.525 0.665 11.99 0.67 ;
      RECT  10.525 0.67 11.995 0.675 ;
      RECT  11.665 0.675 12.0 0.68 ;
      RECT  10.525 0.675 10.755 1.565 ;
      RECT  11.67 0.68 12.005 0.685 ;
      RECT  11.675 0.685 12.01 0.69 ;
      RECT  11.68 0.69 12.015 0.695 ;
      RECT  11.685 0.695 12.02 0.7 ;
      RECT  11.69 0.7 12.025 0.705 ;
      RECT  11.695 0.705 12.03 0.71 ;
      RECT  11.7 0.71 12.035 0.715 ;
      RECT  11.705 0.715 12.04 0.72 ;
      RECT  11.71 0.72 12.045 0.725 ;
      RECT  11.715 0.725 12.05 0.73 ;
      RECT  11.72 0.73 12.055 0.735 ;
      RECT  11.725 0.735 12.06 0.74 ;
      RECT  11.73 0.74 12.065 0.745 ;
      RECT  11.735 0.745 12.07 0.75 ;
      RECT  11.74 0.75 12.94 0.755 ;
      RECT  11.745 0.755 12.94 0.76 ;
      RECT  11.75 0.76 12.94 0.765 ;
      RECT  11.755 0.765 12.94 0.77 ;
      RECT  11.76 0.77 12.94 0.775 ;
      RECT  11.765 0.775 12.94 0.78 ;
      RECT  11.77 0.78 12.94 0.785 ;
      RECT  11.775 0.785 12.94 0.79 ;
      RECT  11.78 0.79 12.94 0.795 ;
      RECT  11.785 0.795 12.94 0.8 ;
      RECT  11.79 0.8 12.94 0.805 ;
      RECT  11.795 0.805 12.94 0.81 ;
      RECT  11.8 0.81 12.94 0.815 ;
      RECT  11.805 0.815 12.94 0.82 ;
      RECT  11.81 0.82 12.94 0.825 ;
      RECT  11.815 0.825 12.94 0.83 ;
      RECT  11.82 0.83 12.94 0.835 ;
      RECT  11.825 0.835 12.94 0.84 ;
      RECT  11.83 0.84 12.94 0.845 ;
      RECT  11.835 0.845 12.94 0.85 ;
      RECT  11.84 0.85 12.94 0.855 ;
      RECT  11.845 0.855 12.94 0.86 ;
      RECT  11.85 0.86 12.94 0.865 ;
      RECT  11.855 0.865 12.94 0.87 ;
      RECT  11.86 0.87 12.94 0.875 ;
      RECT  11.865 0.875 12.94 0.88 ;
      RECT  11.87 0.88 12.94 0.885 ;
      RECT  11.875 0.885 12.94 0.89 ;
      RECT  11.88 0.89 12.94 0.895 ;
      RECT  11.885 0.895 12.94 0.9 ;
      RECT  11.89 0.9 12.94 0.905 ;
      RECT  11.895 0.905 12.94 0.91 ;
      RECT  11.9 0.91 12.94 0.915 ;
      RECT  11.905 0.915 12.94 0.92 ;
      RECT  11.91 0.92 12.94 0.925 ;
      RECT  11.915 0.925 12.94 0.93 ;
      RECT  11.92 0.93 12.94 0.935 ;
      RECT  11.925 0.935 12.94 0.94 ;
      RECT  11.93 0.94 12.94 0.945 ;
      RECT  11.935 0.945 12.94 0.95 ;
      RECT  11.94 0.95 12.94 0.955 ;
      RECT  11.945 0.955 12.94 0.96 ;
      RECT  11.95 0.96 12.94 0.965 ;
      RECT  11.955 0.965 12.94 0.97 ;
      RECT  11.96 0.97 12.94 0.975 ;
      RECT  11.965 0.975 12.94 0.98 ;
      RECT  12.71 0.98 12.94 1.005 ;
      RECT  12.71 1.005 28.945 1.235 ;
      RECT  9.14 1.565 10.755 1.665 ;
      RECT  9.14 1.665 11.315 1.795 ;
      RECT  10.525 1.795 11.315 1.895 ;
      RECT  11.085 1.895 11.315 3.245 ;
      RECT  9.14 3.245 11.315 3.475 ;
      RECT  0.95 0.445 2.615 0.675 ;
      RECT  2.385 0.675 2.615 1.005 ;
      RECT  2.385 1.005 10.25 1.235 ;
      RECT  3.96 1.565 4.3 1.67 ;
      RECT  3.96 1.67 4.305 1.675 ;
      RECT  3.96 1.675 4.31 1.68 ;
      RECT  3.96 1.68 4.315 1.685 ;
      RECT  3.96 1.685 4.32 1.69 ;
      RECT  3.96 1.69 4.325 1.695 ;
      RECT  3.96 1.695 4.33 1.7 ;
      RECT  3.96 1.7 4.335 1.705 ;
      RECT  3.96 1.705 4.34 1.71 ;
      RECT  3.96 1.71 4.345 1.715 ;
      RECT  3.96 1.715 4.35 1.72 ;
      RECT  3.96 1.72 4.355 1.725 ;
      RECT  3.96 1.725 4.36 1.73 ;
      RECT  3.96 1.73 4.365 1.735 ;
      RECT  3.96 1.735 4.37 1.74 ;
      RECT  3.96 1.74 4.375 1.745 ;
      RECT  3.96 1.745 4.38 1.75 ;
      RECT  3.96 1.75 4.385 1.755 ;
      RECT  3.96 1.755 4.39 1.76 ;
      RECT  3.96 1.76 4.395 1.765 ;
      RECT  3.96 1.765 4.4 1.77 ;
      RECT  3.96 1.77 4.405 1.775 ;
      RECT  3.96 1.775 4.41 1.78 ;
      RECT  3.96 1.78 4.415 1.785 ;
      RECT  3.96 1.785 4.42 1.79 ;
      RECT  3.96 1.79 4.425 1.795 ;
      RECT  4.095 1.795 4.43 1.8 ;
      RECT  4.1 1.8 4.435 1.805 ;
      RECT  4.105 1.805 4.44 1.81 ;
      RECT  4.11 1.81 4.445 1.815 ;
      RECT  4.115 1.815 4.45 1.82 ;
      RECT  4.12 1.82 4.455 1.825 ;
      RECT  4.125 1.825 4.46 1.83 ;
      RECT  4.13 1.83 4.465 1.835 ;
      RECT  4.135 1.835 4.47 1.84 ;
      RECT  4.14 1.84 4.475 1.845 ;
      RECT  4.145 1.845 4.48 1.85 ;
      RECT  4.15 1.85 4.485 1.855 ;
      RECT  4.155 1.855 4.49 1.86 ;
      RECT  4.16 1.86 4.495 1.865 ;
      RECT  4.165 1.865 4.5 1.87 ;
      RECT  4.17 1.87 4.505 1.875 ;
      RECT  4.175 1.875 4.51 1.88 ;
      RECT  4.18 1.88 4.515 1.885 ;
      RECT  4.185 1.885 4.52 1.89 ;
      RECT  4.19 1.89 4.525 1.895 ;
      RECT  4.195 1.895 4.53 1.9 ;
      RECT  4.2 1.9 4.535 1.905 ;
      RECT  4.205 1.905 4.54 1.91 ;
      RECT  4.21 1.91 4.545 1.915 ;
      RECT  4.215 1.915 4.55 1.92 ;
      RECT  4.22 1.92 4.555 1.925 ;
      RECT  4.225 1.925 4.56 1.93 ;
      RECT  4.23 1.93 4.565 1.935 ;
      RECT  4.235 1.935 4.57 1.94 ;
      RECT  4.24 1.94 4.575 1.945 ;
      RECT  4.245 1.945 4.58 1.95 ;
      RECT  4.25 1.95 4.585 1.955 ;
      RECT  4.255 1.955 4.59 1.96 ;
      RECT  4.26 1.96 4.595 1.965 ;
      RECT  4.265 1.965 4.595 1.97 ;
      RECT  4.27 1.97 4.595 1.975 ;
      RECT  4.275 1.975 4.595 1.98 ;
      RECT  4.28 1.98 4.595 1.985 ;
      RECT  4.285 1.985 4.595 1.99 ;
      RECT  4.29 1.99 4.595 1.995 ;
      RECT  4.295 1.995 4.595 2.0 ;
      RECT  4.3 2.0 4.595 2.005 ;
      RECT  4.305 2.005 4.595 2.01 ;
      RECT  4.31 2.01 4.595 2.015 ;
      RECT  4.315 2.015 4.595 2.02 ;
      RECT  4.32 2.02 4.595 2.025 ;
      RECT  4.325 2.025 4.595 2.03 ;
      RECT  4.33 2.03 4.595 2.035 ;
      RECT  4.335 2.035 4.595 2.04 ;
      RECT  4.34 2.04 4.595 2.045 ;
      RECT  4.345 2.045 4.595 2.05 ;
      RECT  4.35 2.05 4.595 2.055 ;
      RECT  4.355 2.055 4.595 2.06 ;
      RECT  4.36 2.06 4.595 2.065 ;
      RECT  4.365 2.065 4.595 2.405 ;
      RECT  4.365 2.405 6.33 2.635 ;
      RECT  4.365 2.635 4.595 3.245 ;
      RECT  3.96 3.245 4.595 3.475 ;
      RECT  11.645 2.35 27.61 2.58 ;
      RECT  11.645 2.58 11.875 3.805 ;
      RECT  4.66 1.465 5.715 1.565 ;
      RECT  4.66 1.565 8.785 1.695 ;
      RECT  6.605 1.56 6.835 1.565 ;
      RECT  5.485 1.695 8.785 1.795 ;
      RECT  5.485 1.795 5.715 1.8 ;
      RECT  6.605 1.795 6.835 3.25 ;
      RECT  6.605 3.25 7.395 3.48 ;
      RECT  7.165 3.48 7.395 3.805 ;
      RECT  7.165 3.805 11.875 4.035 ;
      RECT  4.66 3.805 6.835 4.035 ;
      RECT  6.605 4.035 6.835 4.365 ;
      RECT  6.605 4.365 8.78 4.595 ;
      RECT  9.14 4.365 11.02 4.595 ;
      RECT  9.14 4.595 9.37 4.925 ;
      RECT  2.39 4.365 6.275 4.595 ;
      RECT  2.39 4.595 2.62 4.925 ;
      RECT  6.045 4.595 6.275 4.925 ;
      RECT  0.95 4.925 2.62 5.155 ;
      RECT  6.045 4.925 9.37 5.155 ;
  END
END MDN_BUFTS_8
#-----------------------------------------------------------------------
#      Cell        : MDN_BUSH_1
#      Description : Bus holder
#      Equation    : X=keeper(X)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_BUSH_1
  CLASS CORE ;
  FOREIGN MDN_BUSH_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 5.46 11.37 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 -0.14 11.37 0.14 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION INOUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.39 0.37 0.73 0.6 ;
      RECT  0.445 0.6 0.675 1.005 ;
      RECT  0.445 1.005 11.02 1.235 ;
      RECT  9.965 1.235 10.195 3.53 ;
    END
    ANTENNADIFFAREA 2.086 ;
    ANTENNAGATEAREA 0.567 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  9.35 0.37 10.81 0.6 ;
      RECT  1.72 1.565 2.76 1.795 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  8.44 1.565 9.48 1.795 ;
      RECT  0.18 1.565 0.675 1.8 ;
      RECT  0.445 1.8 0.675 2.405 ;
      RECT  0.445 2.405 9.545 2.635 ;
      RECT  0.445 2.635 0.675 3.245 ;
      RECT  0.18 3.245 0.675 3.475 ;
      RECT  1.72 3.245 2.76 3.475 ;
      RECT  3.96 3.245 5.0 3.475 ;
      RECT  6.2 3.245 7.24 3.475 ;
      RECT  8.44 3.245 9.48 3.475 ;
  END
END MDN_BUSH_1
#-----------------------------------------------------------------------
#      Cell        : MDN_CKGTPLS_1
#      Description : Clock Gater, positive clock, synchronous enable, post control
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN):Q=CK&(iq|SE)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_CKGTPLS_1
  CLASS CORE ;
  FOREIGN MDN_CKGTPLS_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 4.365 11.9 5.0 ;
      RECT  10.47 5.0 11.93 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.765 1.565 13.26 1.795 ;
      RECT  12.765 1.795 12.995 3.245 ;
      RECT  12.765 3.245 13.26 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 8.54 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.365 11.02 4.595 ;
      RECT  9.965 4.595 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  4.48 5.46 5.715 5.74 ;
      RECT  1.005 4.925 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  8.96 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 1.005 ;
      RECT  9.14 1.005 10.195 1.235 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.245 1.005 6.22 1.235 ;
      RECT  3.245 1.235 3.475 3.315 ;
      RECT  8.285 0.37 9.69 0.6 ;
      RECT  8.285 0.6 8.515 1.005 ;
      RECT  7.165 1.005 8.515 1.235 ;
      RECT  7.165 1.235 7.395 1.565 ;
      RECT  6.9 1.565 7.395 1.795 ;
      RECT  7.165 1.795 7.395 3.245 ;
      RECT  6.9 3.245 7.395 3.475 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  10.525 1.005 12.94 1.235 ;
      RECT  10.525 1.235 10.755 3.245 ;
      RECT  9.91 3.245 10.755 3.475 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  1.72 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
      RECT  2.685 3.475 2.915 3.545 ;
      RECT  2.685 3.545 4.035 3.775 ;
      RECT  3.805 2.335 4.035 3.545 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 2.405 ;
      RECT  4.87 2.405 6.275 2.635 ;
      RECT  6.045 2.635 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
      RECT  8.44 1.565 10.25 1.795 ;
      RECT  11.085 1.565 11.72 1.795 ;
      RECT  11.085 1.795 11.315 3.245 ;
      RECT  11.085 3.245 11.72 3.475 ;
      RECT  11.085 3.475 11.315 3.805 ;
      RECT  9.405 3.805 11.315 4.035 ;
      RECT  9.405 4.035 9.635 4.365 ;
      RECT  4.925 4.365 9.635 4.595 ;
      RECT  4.925 4.595 5.155 5.0 ;
      RECT  1.51 5.0 5.155 5.23 ;
      RECT  4.365 3.245 5.0 3.475 ;
      RECT  4.365 3.475 4.595 4.005 ;
      RECT  2.38 4.005 4.595 4.235 ;
      RECT  8.845 3.245 9.48 3.475 ;
      RECT  8.845 3.475 9.075 3.805 ;
      RECT  8.44 3.805 9.075 4.035 ;
      RECT  0.14 4.465 4.3 4.695 ;
  END
END MDN_CKGTPLS_1
#-----------------------------------------------------------------------
#      Cell        : MDN_CKGTPLS_2
#      Description : Clock Gater, positive clock, synchronous enable, post control
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN):Q=CK&(iq|SE)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_CKGTPLS_2
  CLASS CORE ;
  FOREIGN MDN_CKGTPLS_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 4.365 11.9 5.0 ;
      RECT  10.47 5.0 11.93 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.92 1.565 13.96 1.795 ;
      RECT  13.325 1.795 13.555 3.245 ;
      RECT  12.92 3.245 13.96 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 8.54 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  9.965 4.365 11.02 4.595 ;
      RECT  9.965 4.595 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  8.96 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 1.005 ;
      RECT  9.14 1.005 10.195 1.235 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.245 1.005 6.22 1.235 ;
      RECT  3.245 1.235 3.475 3.315 ;
      RECT  8.285 0.37 9.69 0.6 ;
      RECT  8.285 0.6 8.515 1.005 ;
      RECT  7.165 1.005 8.515 1.235 ;
      RECT  7.165 1.235 7.395 1.565 ;
      RECT  6.9 1.565 7.395 1.795 ;
      RECT  7.165 1.795 7.395 3.245 ;
      RECT  6.9 3.245 7.395 3.475 ;
      RECT  12.71 0.37 14.17 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  10.525 1.005 12.94 1.235 ;
      RECT  10.525 1.235 10.755 3.245 ;
      RECT  9.91 3.245 10.755 3.475 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
      RECT  2.685 3.475 2.915 3.545 ;
      RECT  2.685 3.545 4.035 3.775 ;
      RECT  3.805 2.35 4.035 3.545 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 2.405 ;
      RECT  4.87 2.405 6.275 2.635 ;
      RECT  6.045 2.635 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
      RECT  8.44 1.565 10.25 1.795 ;
      RECT  11.085 1.565 11.72 1.795 ;
      RECT  11.085 1.795 11.315 3.245 ;
      RECT  11.085 3.245 11.72 3.475 ;
      RECT  11.085 3.475 11.315 3.805 ;
      RECT  9.405 3.805 11.315 4.035 ;
      RECT  9.405 4.035 9.635 4.365 ;
      RECT  4.925 4.365 9.635 4.595 ;
      RECT  4.925 4.595 5.155 5.0 ;
      RECT  1.51 5.0 5.155 5.23 ;
      RECT  4.365 3.245 5.0 3.475 ;
      RECT  4.365 3.475 4.595 4.005 ;
      RECT  2.42 4.005 4.595 4.235 ;
      RECT  8.845 3.245 9.48 3.475 ;
      RECT  8.845 3.475 9.075 3.805 ;
      RECT  8.44 3.805 9.075 4.035 ;
      RECT  0.18 4.465 4.3 4.695 ;
  END
END MDN_CKGTPLS_2
#-----------------------------------------------------------------------
#      Cell        : MDN_CKGTPLS_3
#      Description : Clock Gater, positive clock, synchronous enable, post control
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN):Q=CK&(iq|SE)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_CKGTPLS_3
  CLASS CORE ;
  FOREIGN MDN_CKGTPLS_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 4.365 11.9 5.0 ;
      RECT  10.47 5.0 11.93 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.92 1.565 15.5 1.795 ;
      RECT  14.445 1.795 14.675 3.245 ;
      RECT  12.92 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 4.536 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 8.54 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  9.965 4.365 11.02 4.595 ;
      RECT  9.965 4.595 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  4.48 5.46 5.715 5.74 ;
      RECT  1.005 4.925 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  8.96 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 1.005 ;
      RECT  9.14 1.005 10.195 1.235 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.245 1.005 6.22 1.235 ;
      RECT  3.245 1.235 3.475 3.315 ;
      RECT  8.285 0.37 9.69 0.6 ;
      RECT  8.285 0.6 8.515 1.005 ;
      RECT  7.165 1.005 8.515 1.235 ;
      RECT  7.165 1.235 7.395 1.565 ;
      RECT  6.9 1.565 7.395 1.795 ;
      RECT  7.165 1.795 7.395 3.245 ;
      RECT  6.9 3.245 7.395 3.475 ;
      RECT  14.95 0.37 15.29 0.6 ;
      RECT  14.95 0.6 15.18 1.005 ;
      RECT  12.71 0.37 14.17 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  13.94 0.6 14.17 1.005 ;
      RECT  10.525 1.005 12.94 1.235 ;
      RECT  13.94 1.005 15.18 1.235 ;
      RECT  10.525 1.235 10.755 3.245 ;
      RECT  9.91 3.245 10.755 3.475 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  1.72 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 3.245 ;
      RECT  1.72 3.245 2.355 3.475 ;
      RECT  2.125 3.475 2.355 3.545 ;
      RECT  2.125 3.545 4.035 3.775 ;
      RECT  3.805 2.35 4.035 3.545 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 2.405 ;
      RECT  4.87 2.405 6.275 2.635 ;
      RECT  6.045 2.635 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
      RECT  8.39 1.565 10.25 1.795 ;
      RECT  11.085 1.565 11.72 1.795 ;
      RECT  11.085 1.795 11.315 3.245 ;
      RECT  11.085 3.245 11.72 3.475 ;
      RECT  11.085 3.475 11.315 3.805 ;
      RECT  9.405 3.805 11.315 4.035 ;
      RECT  9.405 4.035 9.635 4.365 ;
      RECT  4.925 4.365 9.635 4.595 ;
      RECT  4.925 4.595 5.155 5.0 ;
      RECT  1.51 5.0 5.155 5.23 ;
      RECT  8.845 3.245 9.48 3.475 ;
      RECT  8.845 3.475 9.075 3.805 ;
      RECT  8.44 3.805 9.075 4.035 ;
      RECT  4.365 3.805 5.0 4.005 ;
      RECT  2.38 4.005 5.0 4.035 ;
      RECT  2.38 4.035 4.595 4.235 ;
      RECT  0.14 4.465 4.3 4.695 ;
  END
END MDN_CKGTPLS_3
#-----------------------------------------------------------------------
#      Cell        : MDN_CKGTPLS_4
#      Description : Clock Gater, positive clock, synchronous enable, post control
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN):Q=CK&(iq|SE)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_CKGTPLS_4
  CLASS CORE ;
  FOREIGN MDN_CKGTPLS_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 4.365 11.9 5.0 ;
      RECT  10.47 5.0 11.93 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.92 1.565 16.2 1.795 ;
      RECT  14.445 1.795 14.675 3.245 ;
      RECT  12.92 3.245 16.2 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 8.54 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.925 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  9.965 4.365 11.02 4.595 ;
      RECT  9.965 4.595 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  4.48 5.46 5.715 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.695 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  8.96 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 1.005 ;
      RECT  9.14 1.005 10.195 1.235 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.245 1.005 6.22 1.235 ;
      RECT  3.245 1.235 3.475 3.315 ;
      RECT  8.285 0.37 9.69 0.6 ;
      RECT  8.285 0.6 8.515 1.005 ;
      RECT  7.165 1.005 8.515 1.235 ;
      RECT  7.165 1.235 7.395 1.565 ;
      RECT  6.9 1.565 7.395 1.795 ;
      RECT  7.165 1.795 7.395 3.245 ;
      RECT  6.9 3.245 7.395 3.475 ;
      RECT  14.95 0.37 16.41 0.6 ;
      RECT  14.95 0.6 15.18 1.005 ;
      RECT  12.71 0.37 14.17 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  13.94 0.6 14.17 1.005 ;
      RECT  10.525 1.005 12.94 1.235 ;
      RECT  13.94 1.005 15.18 1.235 ;
      RECT  10.525 1.235 10.755 3.245 ;
      RECT  9.91 3.245 10.755 3.475 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
      RECT  2.685 3.475 2.915 3.545 ;
      RECT  2.685 3.545 4.035 3.775 ;
      RECT  3.805 2.35 4.035 3.545 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 2.405 ;
      RECT  4.87 2.405 6.275 2.635 ;
      RECT  6.045 2.635 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
      RECT  8.44 1.565 10.25 1.795 ;
      RECT  11.085 1.565 11.72 1.795 ;
      RECT  11.085 1.795 11.315 3.245 ;
      RECT  11.085 3.245 11.72 3.475 ;
      RECT  11.085 3.475 11.315 3.805 ;
      RECT  9.405 3.805 11.315 4.035 ;
      RECT  9.405 4.035 9.635 4.365 ;
      RECT  4.925 4.365 9.635 4.595 ;
      RECT  4.925 4.595 5.155 5.0 ;
      RECT  1.51 5.0 5.155 5.23 ;
      RECT  8.845 3.245 9.48 3.475 ;
      RECT  8.845 3.475 9.075 3.805 ;
      RECT  8.44 3.805 9.075 4.035 ;
      RECT  4.365 3.805 5.0 4.005 ;
      RECT  2.38 4.005 5.0 4.035 ;
      RECT  2.38 4.035 4.595 4.235 ;
      RECT  0.18 4.465 4.3 4.695 ;
  END
END MDN_CKGTPLS_4
#-----------------------------------------------------------------------
#      Cell        : MDN_CKGTPLS_6
#      Description : Clock Gater, positive clock, synchronous enable, post control
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN):Q=CK&(iq|SE)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_CKGTPLS_6
  CLASS CORE ;
  FOREIGN MDN_CKGTPLS_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 24.64 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.885 4.365 15.235 4.595 ;
      RECT  13.885 4.595 14.115 5.0 ;
      RECT  15.005 4.595 15.235 5.0 ;
      RECT  13.83 5.0 14.17 5.23 ;
      RECT  14.95 5.0 16.41 5.23 ;
      RECT  16.1 4.365 16.38 5.0 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.4 1.565 22.92 1.795 ;
      RECT  20.045 1.795 20.275 3.245 ;
      RECT  17.4 3.245 22.92 3.475 ;
    END
    ANTENNADIFFAREA 9.072 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 10.78 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.81 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 21.84 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  14.445 4.905 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 24.64 5.74 ;
      LAYER VIA12 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  24.23 5.47 24.49 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 -0.14 24.81 0.14 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  18.925 -0.14 21.395 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  11.76 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  6.045 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  6.045 0.14 6.275 0.89 ;
      RECT  6.045 0.89 6.54 1.12 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 24.64 0.14 ;
      LAYER VIA12 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  20.31 -0.13 20.57 0.13 ;
      RECT  20.87 -0.13 21.13 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  8.22 0.37 8.57 0.6 ;
      RECT  8.22 0.6 8.45 1.005 ;
      RECT  7.11 0.37 7.45 0.6 ;
      RECT  7.22 0.6 7.45 1.005 ;
      RECT  7.22 1.005 8.45 1.235 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  11.59 0.37 11.93 0.6 ;
      RECT  11.7 0.6 11.93 1.005 ;
      RECT  8.68 1.005 12.94 1.235 ;
      RECT  8.68 1.235 8.91 1.565 ;
      RECT  8.285 1.565 8.91 1.795 ;
      RECT  8.285 1.795 8.515 3.245 ;
      RECT  8.285 3.245 8.78 3.475 ;
      RECT  21.67 0.37 23.13 0.6 ;
      RECT  21.67 0.6 21.9 1.005 ;
      RECT  19.43 0.37 20.89 0.6 ;
      RECT  19.43 0.6 19.66 1.005 ;
      RECT  20.66 0.6 20.89 1.005 ;
      RECT  17.19 0.37 18.65 0.6 ;
      RECT  17.19 0.6 17.42 1.005 ;
      RECT  18.42 0.6 18.65 1.005 ;
      RECT  14.445 1.005 17.42 1.235 ;
      RECT  18.42 1.005 19.66 1.235 ;
      RECT  20.66 1.005 21.9 1.235 ;
      RECT  14.445 1.235 14.675 3.245 ;
      RECT  11.38 3.245 15.5 3.475 ;
      RECT  0.14 1.005 2.76 1.235 ;
      RECT  3.96 1.005 5.77 1.235 ;
      RECT  3.19 1.565 6.275 1.795 ;
      RECT  6.045 1.795 6.275 2.39 ;
      RECT  3.19 1.795 3.42 3.03 ;
      RECT  6.045 2.39 7.225 2.62 ;
      RECT  3.19 3.03 3.53 3.26 ;
      RECT  6.9 1.565 7.955 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  6.9 3.245 7.955 3.475 ;
      RECT  9.14 1.565 13.96 1.795 ;
      RECT  15.86 1.565 16.355 1.795 ;
      RECT  16.125 1.795 16.355 3.805 ;
      RECT  13.325 3.805 16.355 4.035 ;
      RECT  13.325 4.035 13.555 4.365 ;
      RECT  4.925 3.805 7.955 4.035 ;
      RECT  7.725 4.035 7.955 4.365 ;
      RECT  4.925 4.035 5.155 5.0 ;
      RECT  7.725 4.365 13.555 4.595 ;
      RECT  1.51 5.0 5.155 5.23 ;
      RECT  3.75 2.405 5.21 2.635 ;
      RECT  3.805 2.635 4.035 3.49 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
      RECT  2.685 3.475 2.915 3.49 ;
      RECT  2.685 3.49 4.035 3.72 ;
      RECT  4.365 3.245 6.54 3.475 ;
      RECT  4.365 3.475 4.595 3.95 ;
      RECT  2.42 3.95 4.595 4.18 ;
      RECT  9.135 3.805 12.49 4.035 ;
      RECT  6.605 4.365 7.24 4.595 ;
      RECT  6.605 4.595 6.835 5.0 ;
      RECT  5.99 5.0 6.835 5.23 ;
      RECT  0.14 4.41 4.3 4.64 ;
  END
END MDN_CKGTPLS_6
#-----------------------------------------------------------------------
#      Cell        : MDN_CKGTPLS_8
#      Description : Clock Gater, positive clock, synchronous enable, post control
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN):Q=CK&(iq|SE)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_CKGTPLS_8
  CLASS CORE ;
  FOREIGN MDN_CKGTPLS_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 26.88 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.885 4.365 15.235 4.595 ;
      RECT  13.885 4.595 14.115 5.0 ;
      RECT  15.005 4.595 15.235 5.0 ;
      RECT  13.83 5.0 14.17 5.23 ;
      RECT  14.95 5.0 16.41 5.23 ;
      RECT  16.1 4.365 16.38 5.0 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.4 1.565 25.16 1.795 ;
      RECT  24.525 1.795 24.755 3.245 ;
      RECT  17.4 3.245 25.16 3.475 ;
    END
    ANTENNADIFFAREA 12.096 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 10.78 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.645 5.46 27.05 5.74 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.08 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 21.84 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.88 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 26.88 5.74 ;
      LAYER VIA12 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 -0.14 27.05 0.14 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  25.645 0.14 25.875 0.7 ;
      RECT  21.165 -0.14 21.84 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.925 -0.14 19.6 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  6.045 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  6.045 0.14 6.275 0.89 ;
      RECT  6.045 0.89 6.54 1.12 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 26.88 0.14 ;
      LAYER VIA12 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  24.79 -0.13 25.05 0.13 ;
      RECT  25.35 -0.13 25.61 0.13 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  8.22 0.37 8.57 0.6 ;
      RECT  8.22 0.6 8.45 1.005 ;
      RECT  7.11 0.37 7.45 0.6 ;
      RECT  7.22 0.6 7.45 1.005 ;
      RECT  7.22 1.005 8.45 1.235 ;
      RECT  7.725 1.235 7.955 3.49 ;
      RECT  3.19 1.565 5.715 1.795 ;
      RECT  3.19 1.795 3.42 3.03 ;
      RECT  5.485 1.795 5.715 3.49 ;
      RECT  3.19 3.03 3.53 3.26 ;
      RECT  5.485 3.49 7.955 3.72 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  11.59 0.37 11.93 0.6 ;
      RECT  11.7 0.6 11.93 1.005 ;
      RECT  8.68 1.005 12.94 1.235 ;
      RECT  8.68 1.235 8.91 1.565 ;
      RECT  8.285 1.565 8.91 1.795 ;
      RECT  8.285 1.795 8.515 3.805 ;
      RECT  8.285 3.805 8.78 4.035 ;
      RECT  23.91 0.37 25.37 0.6 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.005 5.77 1.235 ;
      RECT  14.445 1.005 16.915 1.235 ;
      RECT  16.685 1.235 16.915 2.405 ;
      RECT  14.445 1.235 14.675 3.245 ;
      RECT  16.685 2.405 24.25 2.635 ;
      RECT  11.38 3.245 15.5 3.475 ;
      RECT  6.605 1.565 7.24 1.795 ;
      RECT  6.605 1.795 6.835 2.405 ;
      RECT  5.99 2.405 6.835 2.635 ;
      RECT  6.605 2.635 6.835 3.03 ;
      RECT  6.605 3.03 7.24 3.26 ;
      RECT  9.14 1.565 13.96 1.795 ;
      RECT  15.86 1.565 16.355 1.795 ;
      RECT  16.125 1.795 16.355 3.805 ;
      RECT  13.325 3.805 16.355 4.035 ;
      RECT  13.325 4.035 13.555 4.365 ;
      RECT  7.165 4.365 13.555 4.41 ;
      RECT  4.925 4.41 13.555 4.595 ;
      RECT  4.925 4.595 7.395 4.64 ;
      RECT  4.925 4.64 5.155 5.0 ;
      RECT  1.51 5.0 5.155 5.23 ;
      RECT  3.805 2.405 5.21 2.635 ;
      RECT  3.805 2.635 4.035 3.49 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
      RECT  2.685 3.475 2.915 3.49 ;
      RECT  2.685 3.49 4.035 3.72 ;
      RECT  9.14 3.805 12.49 4.035 ;
      RECT  2.42 3.95 6.54 4.18 ;
      RECT  0.18 4.42 4.3 4.65 ;
  END
END MDN_CKGTPLS_8
#-----------------------------------------------------------------------
#      Cell        : MDN_CKGTPLT_1
#      Description : Clock Gater, positive clock, synchronous enable, pre control
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN|SE):Q=CK&iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_CKGTPLT_1
  CLASS CORE ;
  FOREIGN MDN_CKGTPLT_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 9.66 2.355 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.765 1.565 13.26 1.795 ;
      RECT  12.765 1.795 12.995 3.245 ;
      RECT  12.765 3.245 13.26 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.14 4.365 12.435 4.595 ;
      RECT  12.205 4.595 12.435 5.46 ;
      RECT  11.76 5.46 13.61 5.74 ;
      RECT  5.485 4.945 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.945 7.955 5.46 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  8.96 -0.14 9.635 0.14 ;
      RECT  9.405 0.14 9.635 1.005 ;
      RECT  9.14 1.005 9.635 1.235 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.6 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.595 0.6 ;
      RECT  4.365 0.6 4.595 0.83 ;
      RECT  4.365 0.83 7.185 1.06 ;
      RECT  6.955 1.06 7.185 1.785 ;
      RECT  6.605 1.785 7.185 2.015 ;
      RECT  6.605 2.015 6.835 3.03 ;
      RECT  6.605 3.03 7.24 3.26 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  9.965 1.005 12.94 1.235 ;
      RECT  9.965 1.235 10.195 3.5 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  7.725 1.005 8.78 1.235 ;
      RECT  7.725 1.235 7.955 2.405 ;
      RECT  7.11 2.405 7.955 2.635 ;
      RECT  7.725 2.635 7.955 3.545 ;
      RECT  2.685 2.35 2.915 3.545 ;
      RECT  2.685 3.545 7.955 3.775 ;
      RECT  7.725 3.775 7.955 3.805 ;
      RECT  7.725 3.805 8.78 4.035 ;
      RECT  3.96 1.29 6.54 1.52 ;
      RECT  10.525 1.565 11.72 1.795 ;
      RECT  10.525 1.795 10.755 3.245 ;
      RECT  10.525 3.245 11.72 3.475 ;
      RECT  4.66 1.75 5.155 1.98 ;
      RECT  4.925 1.98 5.155 2.405 ;
      RECT  4.925 2.405 6.33 2.635 ;
      RECT  4.925 2.635 5.155 3.03 ;
      RECT  4.66 3.03 5.155 3.26 ;
      RECT  3.245 1.51 3.475 3.315 ;
      RECT  2.42 4.005 6.54 4.235 ;
      RECT  1.72 4.465 4.3 4.695 ;
      RECT  4.98 4.485 8.515 4.715 ;
      RECT  4.98 4.715 5.21 5.0 ;
      RECT  8.285 4.715 8.515 5.0 ;
      RECT  3.19 5.0 5.21 5.23 ;
      RECT  8.285 5.0 11.93 5.23 ;
  END
END MDN_CKGTPLT_1
#-----------------------------------------------------------------------
#      Cell        : MDN_CKGTPLT_2
#      Description : Clock Gater, positive clock, synchronous enable, pre control
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN|SE):Q=CK&iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_CKGTPLT_2
  CLASS CORE ;
  FOREIGN MDN_CKGTPLT_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 9.66 2.355 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.92 1.565 13.96 1.795 ;
      RECT  13.325 1.795 13.555 3.245 ;
      RECT  12.92 3.245 13.96 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  9.14 4.365 12.435 4.595 ;
      RECT  12.205 4.595 12.435 5.46 ;
      RECT  11.03 5.46 12.435 5.74 ;
      RECT  7.725 4.945 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.945 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  8.96 -0.14 9.635 0.14 ;
      RECT  9.405 0.14 9.635 1.005 ;
      RECT  9.14 1.005 9.635 1.235 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.6 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.595 0.6 ;
      RECT  4.365 0.6 4.595 0.83 ;
      RECT  4.365 0.83 7.185 1.06 ;
      RECT  6.955 1.06 7.185 1.785 ;
      RECT  6.605 1.785 7.185 2.015 ;
      RECT  6.605 2.015 6.835 3.03 ;
      RECT  6.605 3.03 7.24 3.26 ;
      RECT  12.71 0.37 14.17 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  9.965 1.005 12.94 1.235 ;
      RECT  9.965 1.235 10.195 3.5 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  7.725 1.005 8.78 1.235 ;
      RECT  7.725 1.235 7.955 2.405 ;
      RECT  7.11 2.405 7.955 2.635 ;
      RECT  7.725 2.635 7.955 3.545 ;
      RECT  2.685 2.35 2.915 3.545 ;
      RECT  2.685 3.545 7.955 3.775 ;
      RECT  7.725 3.775 7.955 3.805 ;
      RECT  7.725 3.805 8.78 4.035 ;
      RECT  3.96 1.29 6.54 1.52 ;
      RECT  10.525 1.565 11.72 1.795 ;
      RECT  10.525 1.795 10.755 3.245 ;
      RECT  10.525 3.245 11.72 3.475 ;
      RECT  4.66 1.75 5.155 1.98 ;
      RECT  4.925 1.98 5.155 2.405 ;
      RECT  4.925 2.405 6.33 2.635 ;
      RECT  4.925 2.635 5.155 3.03 ;
      RECT  4.66 3.03 5.155 3.26 ;
      RECT  3.245 1.51 3.475 3.315 ;
      RECT  2.42 4.005 6.54 4.235 ;
      RECT  1.72 4.465 4.3 4.695 ;
      RECT  4.98 4.485 8.515 4.715 ;
      RECT  4.98 4.715 5.21 5.0 ;
      RECT  8.285 4.715 8.515 5.0 ;
      RECT  3.175 5.0 5.21 5.23 ;
      RECT  8.285 5.0 11.93 5.23 ;
  END
END MDN_CKGTPLT_2
#-----------------------------------------------------------------------
#      Cell        : MDN_CKGTPLT_3
#      Description : Clock Gater, positive clock, synchronous enable, pre control
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN|SE):Q=CK&iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_CKGTPLT_3
  CLASS CORE ;
  FOREIGN MDN_CKGTPLT_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 9.66 2.355 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.92 1.565 15.5 1.795 ;
      RECT  13.325 1.795 13.555 3.245 ;
      RECT  12.92 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 4.536 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  9.14 4.365 12.435 4.595 ;
      RECT  12.205 4.595 12.435 5.46 ;
      RECT  11.03 5.46 12.435 5.74 ;
      RECT  7.725 4.945 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.945 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  8.96 -0.14 9.635 0.14 ;
      RECT  9.405 0.14 9.635 1.005 ;
      RECT  9.14 1.005 9.635 1.235 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.6 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.595 0.6 ;
      RECT  4.365 0.6 4.595 0.83 ;
      RECT  4.365 0.83 7.185 1.06 ;
      RECT  6.955 1.06 7.185 1.785 ;
      RECT  6.605 1.785 7.185 2.015 ;
      RECT  6.605 2.015 6.835 3.03 ;
      RECT  6.605 3.03 7.24 3.26 ;
      RECT  12.71 0.37 14.17 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  9.965 1.005 12.94 1.235 ;
      RECT  9.965 1.235 10.195 3.49 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  7.725 1.005 8.78 1.235 ;
      RECT  7.725 1.235 7.955 2.405 ;
      RECT  7.11 2.405 7.955 2.635 ;
      RECT  7.725 2.635 7.955 3.545 ;
      RECT  2.685 2.35 2.915 3.545 ;
      RECT  2.685 3.545 7.955 3.775 ;
      RECT  7.725 3.775 7.955 3.805 ;
      RECT  7.725 3.805 8.78 4.035 ;
      RECT  3.96 1.29 6.54 1.52 ;
      RECT  10.525 1.565 11.72 1.795 ;
      RECT  10.525 1.795 10.755 3.245 ;
      RECT  10.525 3.245 11.72 3.475 ;
      RECT  4.66 1.75 5.155 1.98 ;
      RECT  4.925 1.98 5.155 2.405 ;
      RECT  4.925 2.405 6.33 2.635 ;
      RECT  4.925 2.635 5.155 3.03 ;
      RECT  4.66 3.03 5.155 3.26 ;
      RECT  13.945 2.405 15.29 2.635 ;
      RECT  3.245 1.51 3.475 3.315 ;
      RECT  2.42 4.005 6.54 4.235 ;
      RECT  1.72 4.465 4.3 4.695 ;
      RECT  4.98 4.485 8.515 4.715 ;
      RECT  4.98 4.715 5.21 5.0 ;
      RECT  8.285 4.715 8.515 5.0 ;
      RECT  3.19 5.0 5.21 5.23 ;
      RECT  8.285 5.0 11.93 5.23 ;
  END
END MDN_CKGTPLT_3
#-----------------------------------------------------------------------
#      Cell        : MDN_CKGTPLT_4
#      Description : Clock Gater, positive clock, synchronous enable, pre control
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN|SE):Q=CK&iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_CKGTPLT_4
  CLASS CORE ;
  FOREIGN MDN_CKGTPLT_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 9.66 2.355 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.92 1.565 16.2 1.795 ;
      RECT  13.325 1.795 13.555 3.245 ;
      RECT  12.92 3.245 16.2 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  9.14 4.365 12.435 4.595 ;
      RECT  12.205 4.595 12.435 5.46 ;
      RECT  11.03 5.46 12.435 5.74 ;
      RECT  7.725 4.945 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.945 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  0.18 4.395 0.675 4.625 ;
      RECT  0.445 4.625 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  8.96 -0.14 9.635 0.14 ;
      RECT  9.405 0.14 9.635 1.005 ;
      RECT  9.14 1.005 9.635 1.235 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.6 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.595 0.6 ;
      RECT  4.365 0.6 4.595 0.83 ;
      RECT  4.365 0.83 7.185 1.06 ;
      RECT  6.955 1.06 7.185 1.785 ;
      RECT  6.605 1.785 7.185 2.015 ;
      RECT  6.605 2.015 6.835 3.03 ;
      RECT  6.605 3.03 7.24 3.26 ;
      RECT  12.71 0.37 14.17 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  9.965 1.005 12.94 1.235 ;
      RECT  9.965 1.235 10.195 3.5 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  7.725 1.005 8.78 1.235 ;
      RECT  7.725 1.235 7.955 2.405 ;
      RECT  7.11 2.405 7.955 2.635 ;
      RECT  7.725 2.635 7.955 3.545 ;
      RECT  2.685 2.35 2.915 3.545 ;
      RECT  2.685 3.545 7.955 3.775 ;
      RECT  7.725 3.775 7.955 3.805 ;
      RECT  7.725 3.805 8.78 4.035 ;
      RECT  3.96 1.29 6.54 1.52 ;
      RECT  11.085 1.565 11.72 1.795 ;
      RECT  11.085 1.795 11.315 2.405 ;
      RECT  10.47 2.405 11.315 2.635 ;
      RECT  11.085 2.635 11.315 3.245 ;
      RECT  11.085 3.245 11.72 3.475 ;
      RECT  4.66 1.75 5.155 1.98 ;
      RECT  4.925 1.98 5.155 2.405 ;
      RECT  4.925 2.405 6.33 2.635 ;
      RECT  4.925 2.635 5.155 3.03 ;
      RECT  4.66 3.03 5.155 3.26 ;
      RECT  13.885 2.125 16.355 2.355 ;
      RECT  13.885 2.355 14.115 2.69 ;
      RECT  15.005 2.355 15.235 2.69 ;
      RECT  16.125 2.355 16.355 2.69 ;
      RECT  3.245 1.51 3.475 3.315 ;
      RECT  2.42 4.005 6.54 4.235 ;
      RECT  1.72 4.465 4.3 4.695 ;
      RECT  4.98 4.485 8.515 4.715 ;
      RECT  8.285 4.715 8.515 4.925 ;
      RECT  4.98 4.715 5.21 5.0 ;
      RECT  8.285 4.925 11.93 5.155 ;
      RECT  3.19 5.0 5.21 5.23 ;
      RECT  11.59 5.155 11.93 5.23 ;
  END
END MDN_CKGTPLT_4
#-----------------------------------------------------------------------
#      Cell        : MDN_CKGTPLT_6
#      Description : Clock Gater, positive clock, synchronous enable, pre control
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN|SE):Q=CK&iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_CKGTPLT_6
  CLASS CORE ;
  FOREIGN MDN_CKGTPLT_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 10.78 2.355 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.16 1.565 20.68 1.795 ;
      RECT  20.045 1.795 20.275 3.245 ;
      RECT  15.16 3.245 20.68 3.475 ;
    END
    ANTENNADIFFAREA 9.072 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 22.57 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  9.965 4.945 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.945 12.435 5.46 ;
      RECT  5.485 4.945 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.945 7.955 5.46 ;
      RECT  0.18 4.395 0.675 4.625 ;
      RECT  0.445 4.625 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  20.31 5.47 20.57 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 22.57 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.6 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  20.31 -0.13 20.57 0.13 ;
      RECT  20.87 -0.13 21.13 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.595 0.6 ;
      RECT  4.365 0.6 4.595 0.83 ;
      RECT  4.365 0.83 7.185 1.06 ;
      RECT  6.955 1.06 7.185 1.785 ;
      RECT  6.605 1.785 7.185 2.015 ;
      RECT  6.605 2.015 6.835 3.03 ;
      RECT  6.605 3.03 7.24 3.26 ;
      RECT  11.59 0.37 13.555 0.6 ;
      RECT  13.325 0.6 13.555 1.005 ;
      RECT  13.325 1.005 14.115 1.235 ;
      RECT  13.885 1.235 14.115 3.245 ;
      RECT  13.62 3.245 14.115 3.475 ;
      RECT  19.43 0.37 20.89 0.6 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  7.725 1.005 8.78 1.235 ;
      RECT  7.725 1.235 7.955 2.405 ;
      RECT  7.11 2.405 7.955 2.635 ;
      RECT  7.725 2.635 7.955 3.545 ;
      RECT  2.685 2.35 2.915 3.545 ;
      RECT  2.685 3.545 7.955 3.775 ;
      RECT  7.725 3.775 7.955 3.805 ;
      RECT  7.725 3.805 8.78 4.035 ;
      RECT  9.14 1.005 12.49 1.235 ;
      RECT  3.96 1.29 6.54 1.52 ;
      RECT  4.66 1.75 5.155 1.98 ;
      RECT  4.925 1.98 5.155 2.405 ;
      RECT  4.925 2.405 6.33 2.635 ;
      RECT  4.925 2.635 5.155 3.03 ;
      RECT  4.66 3.03 5.155 3.26 ;
      RECT  15.005 2.35 15.235 2.685 ;
      RECT  14.445 2.685 19.5 2.915 ;
      RECT  16.125 2.35 16.355 2.685 ;
      RECT  17.245 2.35 17.475 2.685 ;
      RECT  18.365 2.35 18.595 2.685 ;
      RECT  19.27 2.35 19.5 2.685 ;
      RECT  14.445 2.915 14.675 3.805 ;
      RECT  11.38 1.565 13.26 1.795 ;
      RECT  12.765 1.795 12.995 3.805 ;
      RECT  9.14 3.805 14.675 4.035 ;
      RECT  3.245 1.51 3.475 3.315 ;
      RECT  2.42 4.005 6.54 4.235 ;
      RECT  1.72 4.465 4.3 4.695 ;
      RECT  4.98 4.485 14.06 4.715 ;
      RECT  4.98 4.715 5.21 5.0 ;
      RECT  13.83 4.715 14.06 5.0 ;
      RECT  3.19 5.0 5.21 5.23 ;
      RECT  13.83 5.0 14.17 5.23 ;
  END
END MDN_CKGTPLT_6
#-----------------------------------------------------------------------
#      Cell        : MDN_CKGTPLT_8
#      Description : Clock Gater, positive clock, synchronous enable, pre control
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN|SE):Q=CK&iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_CKGTPLT_8
  CLASS CORE ;
  FOREIGN MDN_CKGTPLT_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 24.64 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 10.78 2.355 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.16 1.565 22.92 1.795 ;
      RECT  22.285 1.795 22.515 3.245 ;
      RECT  15.16 3.245 22.92 3.475 ;
    END
    ANTENNADIFFAREA 12.096 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 24.81 5.74 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  9.965 4.945 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.945 12.435 5.46 ;
      RECT  5.485 4.945 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.945 7.955 5.46 ;
      RECT  0.18 4.395 0.675 4.625 ;
      RECT  0.445 4.625 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 24.64 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  22.55 5.47 22.81 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  24.23 5.47 24.49 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 24.81 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  18.925 -0.14 19.6 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.6 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 24.64 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  22.55 -0.13 22.81 0.13 ;
      RECT  23.11 -0.13 23.37 0.13 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.595 0.6 ;
      RECT  4.365 0.6 4.595 0.83 ;
      RECT  4.365 0.83 7.185 1.06 ;
      RECT  6.955 1.06 7.185 1.785 ;
      RECT  6.605 1.785 7.185 2.015 ;
      RECT  6.605 2.015 6.835 3.03 ;
      RECT  6.605 3.03 7.24 3.26 ;
      RECT  11.59 0.37 13.555 0.6 ;
      RECT  13.325 0.6 13.555 1.005 ;
      RECT  13.325 1.005 14.115 1.235 ;
      RECT  13.885 1.235 14.115 3.245 ;
      RECT  13.62 3.245 14.115 3.475 ;
      RECT  21.67 0.37 23.13 0.6 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  7.725 1.005 8.78 1.235 ;
      RECT  7.725 1.235 7.955 2.405 ;
      RECT  7.11 2.405 7.955 2.635 ;
      RECT  7.725 2.635 7.955 3.545 ;
      RECT  2.685 2.35 2.915 3.545 ;
      RECT  2.685 3.545 7.955 3.775 ;
      RECT  7.725 3.775 7.955 3.805 ;
      RECT  7.725 3.805 8.78 4.035 ;
      RECT  9.14 1.005 12.49 1.235 ;
      RECT  3.96 1.29 6.54 1.52 ;
      RECT  4.66 1.75 5.155 1.98 ;
      RECT  4.925 1.98 5.155 2.405 ;
      RECT  4.925 2.405 6.33 2.635 ;
      RECT  4.925 2.635 5.155 3.03 ;
      RECT  4.66 3.03 5.155 3.26 ;
      RECT  15.005 2.35 15.235 2.685 ;
      RECT  14.445 2.685 21.955 2.915 ;
      RECT  16.125 2.35 16.355 2.685 ;
      RECT  17.245 2.35 17.475 2.685 ;
      RECT  18.365 2.35 18.595 2.685 ;
      RECT  19.485 2.35 19.715 2.685 ;
      RECT  20.605 2.35 20.835 2.685 ;
      RECT  21.725 2.35 21.955 2.685 ;
      RECT  14.445 2.915 14.675 3.805 ;
      RECT  11.38 1.565 13.26 1.795 ;
      RECT  12.765 1.795 12.995 3.805 ;
      RECT  9.14 3.805 14.675 4.035 ;
      RECT  3.245 1.51 3.475 3.315 ;
      RECT  2.42 4.005 6.54 4.235 ;
      RECT  1.72 4.465 4.3 4.695 ;
      RECT  4.98 4.485 14.06 4.715 ;
      RECT  4.98 4.715 5.21 5.0 ;
      RECT  13.83 4.715 14.06 5.0 ;
      RECT  3.19 5.0 5.21 5.23 ;
      RECT  13.83 5.0 14.17 5.23 ;
  END
END MDN_CKGTPLT_8
#-----------------------------------------------------------------------
#      Cell        : MDN_DEL_R16_1
#      Description : Delay buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_DEL_R16_1
  CLASS CORE ;
  FOREIGN MDN_DEL_R16_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 2.125 11.9 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.1 4.365 18.595 4.595 ;
      RECT  18.365 4.595 18.595 5.46 ;
      RECT  17.92 5.46 18.595 5.74 ;
      RECT  15.86 4.365 16.355 4.595 ;
      RECT  16.125 4.595 16.355 5.46 ;
      RECT  15.68 5.46 16.355 5.74 ;
      RECT  9.14 4.365 9.635 4.595 ;
      RECT  9.405 4.595 9.635 5.46 ;
      RECT  9.405 5.46 12.435 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  6.9 4.365 7.395 4.595 ;
      RECT  7.165 4.595 7.395 5.46 ;
      RECT  6.72 5.46 7.395 5.74 ;
      RECT  4.66 4.365 5.155 4.595 ;
      RECT  4.925 4.595 5.155 5.46 ;
      RECT  4.48 5.46 5.155 5.74 ;
      RECT  2.42 4.365 2.915 4.595 ;
      RECT  2.685 4.595 2.915 5.46 ;
      RECT  2.24 5.46 2.915 5.74 ;
      RECT  -0.17 5.46 0.56 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  18.07 5.47 18.33 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.73 ;
      RECT  16.685 -0.14 18.595 0.14 ;
      RECT  16.685 0.14 16.915 1.005 ;
      RECT  18.365 0.14 18.595 1.005 ;
      RECT  15.82 1.005 16.915 1.235 ;
      RECT  18.1 1.005 18.595 1.235 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.965 0.14 10.195 1.005 ;
      RECT  9.1 1.005 10.195 1.235 ;
      RECT  5.04 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 1.005 ;
      RECT  4.62 1.005 7.255 1.235 ;
      RECT  2.685 -0.14 3.36 0.14 ;
      RECT  2.685 0.14 2.915 1.005 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  18.07 -0.13 18.33 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  21.725 1.565 22.22 1.795 ;
      RECT  21.725 1.795 21.955 3.245 ;
      RECT  21.725 3.245 22.22 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.245 0.37 5.215 0.6 ;
      RECT  3.245 0.6 3.475 1.565 ;
      RECT  2.125 1.565 4.3 1.795 ;
      RECT  2.125 1.795 2.355 2.405 ;
      RECT  3.245 1.795 3.475 3.245 ;
      RECT  0.615 2.405 2.355 2.635 ;
      RECT  3.245 3.245 4.3 3.475 ;
      RECT  5.99 0.37 9.7 0.6 ;
      RECT  7.725 0.6 7.955 1.565 ;
      RECT  7.725 1.565 8.78 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  7.725 3.245 8.78 3.475 ;
      RECT  7.725 3.475 7.955 3.53 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  10.485 1.005 12.94 1.235 ;
      RECT  10.485 1.235 10.715 1.565 ;
      RECT  9.91 1.565 10.715 1.795 ;
      RECT  9.91 1.795 10.14 2.405 ;
      RECT  8.23 2.405 10.14 2.635 ;
      RECT  9.91 2.635 10.14 3.245 ;
      RECT  9.91 3.245 10.25 3.475 ;
      RECT  14.965 0.37 16.42 0.6 ;
      RECT  14.965 0.6 15.195 1.565 ;
      RECT  12.86 1.565 15.5 1.795 ;
      RECT  13.325 1.795 13.555 3.245 ;
      RECT  12.86 3.245 15.5 3.475 ;
      RECT  21.67 0.37 22.01 0.6 ;
      RECT  21.67 0.6 21.9 1.005 ;
      RECT  19.43 0.37 19.77 0.6 ;
      RECT  19.485 0.6 19.715 1.005 ;
      RECT  19.485 1.005 21.9 1.235 ;
      RECT  21.165 1.235 21.395 3.245 ;
      RECT  20.3 3.245 21.395 3.475 ;
      RECT  17.205 1.005 17.74 1.235 ;
      RECT  17.205 1.235 17.435 1.565 ;
      RECT  16.63 1.565 17.435 1.795 ;
      RECT  16.63 1.795 16.86 2.405 ;
      RECT  13.8 2.405 16.86 2.635 ;
      RECT  16.63 2.635 16.86 3.245 ;
      RECT  16.63 3.245 18.595 3.475 ;
      RECT  18.365 2.33 18.595 3.245 ;
      RECT  5.38 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 2.405 ;
      RECT  3.75 2.405 7.24 2.635 ;
      RECT  6.045 2.635 6.275 3.245 ;
      RECT  5.38 3.245 6.54 3.475 ;
      RECT  11.085 1.565 11.72 1.795 ;
      RECT  11.085 1.795 11.315 2.125 ;
      RECT  10.525 2.125 11.315 2.355 ;
      RECT  10.525 2.355 10.755 3.805 ;
      RECT  1.565 1.005 2.06 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  0.13 1.565 1.795 1.795 ;
      RECT  0.13 1.795 0.36 3.245 ;
      RECT  0.13 3.245 2.915 3.475 ;
      RECT  2.685 2.32 2.915 3.245 ;
      RECT  2.685 3.475 2.915 3.805 ;
      RECT  2.685 3.805 11.72 4.035 ;
      RECT  17.805 1.565 19.98 1.795 ;
      RECT  17.805 1.795 18.035 2.405 ;
      RECT  19.485 1.795 19.715 2.405 ;
      RECT  17.19 2.405 18.035 2.635 ;
      RECT  19.485 2.405 20.765 2.635 ;
      RECT  19.485 2.635 19.715 3.245 ;
      RECT  18.825 3.245 19.98 3.475 ;
      RECT  9.91 4.365 11.02 4.595 ;
      RECT  11.645 4.365 13.26 4.595 ;
      RECT  11.645 4.595 11.875 5.0 ;
      RECT  10.47 5.0 11.875 5.23 ;
  END
END MDN_DEL_R16_1
#-----------------------------------------------------------------------
#      Cell        : MDN_DEL_R32_1
#      Description : Delay buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_DEL_R32_1
  CLASS CORE ;
  FOREIGN MDN_DEL_R32_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 29.12 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  28.445 4.365 28.94 4.595 ;
      RECT  28.445 4.595 28.675 5.46 ;
      RECT  28.445 5.46 29.29 5.74 ;
      RECT  25.645 4.87 25.875 5.46 ;
      RECT  25.645 5.46 26.32 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  17.75 5.46 19.155 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 29.12 5.74 ;
      LAYER VIA12 ;
      RECT  28.71 5.47 28.97 5.73 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  18.07 5.47 18.33 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  28.445 -0.14 29.29 0.14 ;
      RECT  28.445 0.14 28.675 1.005 ;
      RECT  28.445 1.005 28.94 1.235 ;
      RECT  25.2 -0.14 25.875 0.14 ;
      RECT  25.645 0.14 25.875 0.73 ;
      RECT  17.75 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  5.485 -0.14 6.89 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 29.12 0.14 ;
      LAYER VIA12 ;
      RECT  28.71 -0.13 28.97 0.13 ;
      RECT  25.35 -0.13 25.61 0.13 ;
      RECT  18.07 -0.13 18.33 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 1.565 26.7 1.795 ;
      RECT  25.645 1.795 25.875 3.245 ;
      RECT  25.645 3.245 26.7 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.83 0.37 5.21 0.6 ;
      RECT  1.83 0.6 2.06 1.565 ;
      RECT  1.005 1.565 2.06 1.795 ;
      RECT  1.005 1.795 1.235 3.245 ;
      RECT  0.95 3.245 2.06 3.475 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  2.315 1.005 6.22 1.235 ;
      RECT  2.315 1.235 2.545 2.405 ;
      RECT  1.51 2.405 2.545 2.635 ;
      RECT  2.315 2.635 2.545 3.245 ;
      RECT  2.315 3.245 3.53 3.475 ;
      RECT  8.535 0.37 11.93 0.6 ;
      RECT  8.535 0.6 8.765 1.565 ;
      RECT  7.725 1.565 8.78 1.795 ;
      RECT  7.725 1.795 7.955 2.405 ;
      RECT  2.795 2.405 7.955 2.635 ;
      RECT  7.725 2.635 7.955 3.245 ;
      RECT  7.725 3.245 8.78 3.475 ;
      RECT  12.71 0.37 14.17 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  9.035 1.005 12.94 1.235 ;
      RECT  9.035 1.235 9.265 2.405 ;
      RECT  8.23 2.405 9.265 2.635 ;
      RECT  9.035 2.635 9.265 3.245 ;
      RECT  9.035 3.245 10.2 3.475 ;
      RECT  15.27 0.37 18.65 0.6 ;
      RECT  15.27 0.6 15.5 1.565 ;
      RECT  14.445 1.565 15.5 1.795 ;
      RECT  14.445 1.795 14.675 2.405 ;
      RECT  9.515 2.405 14.675 2.635 ;
      RECT  14.445 2.635 14.675 3.245 ;
      RECT  14.445 3.245 15.5 3.475 ;
      RECT  19.43 0.37 20.895 0.6 ;
      RECT  19.43 0.6 19.66 1.005 ;
      RECT  15.755 1.005 19.66 1.235 ;
      RECT  15.755 1.235 15.985 2.405 ;
      RECT  14.95 2.405 15.985 2.635 ;
      RECT  15.755 2.635 15.985 3.245 ;
      RECT  15.755 3.245 16.92 3.475 ;
      RECT  21.99 0.37 25.37 0.6 ;
      RECT  21.99 0.6 22.22 1.565 ;
      RECT  21.165 1.565 22.22 1.795 ;
      RECT  21.165 1.795 21.395 2.375 ;
      RECT  16.215 2.375 21.395 2.605 ;
      RECT  21.165 2.605 21.395 3.245 ;
      RECT  21.165 3.245 22.22 3.475 ;
      RECT  27.27 0.37 27.61 0.6 ;
      RECT  27.27 0.6 27.5 1.005 ;
      RECT  22.54 1.005 28.115 1.235 ;
      RECT  22.54 1.235 22.77 2.405 ;
      RECT  27.885 1.235 28.115 2.405 ;
      RECT  21.67 2.405 22.77 2.635 ;
      RECT  27.885 2.405 28.635 2.635 ;
      RECT  22.54 2.635 22.77 3.245 ;
      RECT  22.54 3.245 23.64 3.475 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  6.185 1.565 7.24 1.795 ;
      RECT  10.67 1.565 11.72 1.795 ;
      RECT  12.92 1.565 13.96 1.795 ;
      RECT  17.4 1.565 18.44 1.795 ;
      RECT  19.625 1.565 20.68 1.795 ;
      RECT  24.12 1.565 25.16 1.795 ;
      RECT  27.115 1.51 27.345 2.405 ;
      RECT  26.15 2.405 27.345 2.635 ;
      RECT  27.115 2.635 27.345 3.455 ;
      RECT  3.96 3.245 5.0 3.475 ;
      RECT  6.165 3.245 7.24 3.475 ;
      RECT  10.68 3.245 11.72 3.475 ;
      RECT  12.885 3.245 13.96 3.475 ;
      RECT  17.4 3.245 18.44 3.475 ;
      RECT  19.64 3.245 20.68 3.475 ;
      RECT  24.12 3.245 25.16 3.475 ;
      RECT  25.085 4.365 26.335 4.595 ;
      RECT  25.085 4.595 25.315 5.0 ;
      RECT  26.105 4.595 26.335 5.0 ;
      RECT  22.79 5.0 25.315 5.23 ;
      RECT  26.105 5.0 26.49 5.23 ;
  END
END MDN_DEL_R32_1
#-----------------------------------------------------------------------
#      Cell        : MDN_DEL_R64_1
#      Description : Delay buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_DEL_R64_1
  CLASS CORE ;
  FOREIGN MDN_DEL_R64_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 56 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  55.325 4.365 55.82 4.595 ;
      RECT  55.325 4.595 55.555 5.46 ;
      RECT  55.325 5.46 56.17 5.74 ;
      RECT  52.525 4.87 52.755 5.46 ;
      RECT  52.525 5.46 53.2 5.74 ;
      RECT  45.805 4.9 46.035 5.46 ;
      RECT  44.63 5.46 46.035 5.74 ;
      RECT  39.085 4.9 39.315 5.46 ;
      RECT  38.64 5.46 39.315 5.74 ;
      RECT  32.365 4.9 32.595 5.46 ;
      RECT  32.365 5.46 33.77 5.74 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.645 5.46 27.05 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  17.75 5.46 19.155 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 56.0 5.74 ;
      LAYER VIA12 ;
      RECT  55.59 5.47 55.85 5.73 ;
      RECT  52.79 5.47 53.05 5.73 ;
      RECT  44.95 5.47 45.21 5.73 ;
      RECT  45.51 5.47 45.77 5.73 ;
      RECT  38.79 5.47 39.05 5.73 ;
      RECT  32.63 5.47 32.89 5.73 ;
      RECT  33.19 5.47 33.45 5.73 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  18.07 5.47 18.33 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  55.325 -0.14 56.17 0.14 ;
      RECT  55.325 0.14 55.555 1.005 ;
      RECT  55.325 1.005 55.82 1.235 ;
      RECT  52.525 -0.14 53.2 0.14 ;
      RECT  52.525 0.14 52.755 0.73 ;
      RECT  44.63 -0.14 46.035 0.14 ;
      RECT  45.805 0.14 46.035 0.73 ;
      RECT  38.64 -0.14 39.315 0.14 ;
      RECT  39.085 0.14 39.315 0.73 ;
      RECT  32.365 -0.14 33.77 0.14 ;
      RECT  32.365 0.14 32.595 0.73 ;
      RECT  25.645 -0.14 27.05 0.14 ;
      RECT  25.645 0.14 25.875 0.73 ;
      RECT  17.75 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  5.485 -0.14 6.89 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 56.0 0.14 ;
      LAYER VIA12 ;
      RECT  55.59 -0.13 55.85 0.13 ;
      RECT  52.79 -0.13 53.05 0.13 ;
      RECT  44.95 -0.13 45.21 0.13 ;
      RECT  45.51 -0.13 45.77 0.13 ;
      RECT  38.79 -0.13 39.05 0.13 ;
      RECT  32.63 -0.13 32.89 0.13 ;
      RECT  33.19 -0.13 33.45 0.13 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  18.07 -0.13 18.33 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  52.525 1.565 53.58 1.795 ;
      RECT  52.525 1.795 52.755 3.245 ;
      RECT  52.525 3.245 53.58 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.83 0.37 5.21 0.6 ;
      RECT  1.83 0.6 2.06 1.565 ;
      RECT  1.005 1.565 2.06 1.795 ;
      RECT  1.005 1.795 1.235 3.245 ;
      RECT  1.005 3.245 2.06 3.475 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.25 1.005 6.22 1.235 ;
      RECT  3.25 1.235 3.48 1.565 ;
      RECT  2.315 1.565 3.48 1.795 ;
      RECT  2.315 1.795 2.545 2.405 ;
      RECT  1.51 2.405 2.545 2.635 ;
      RECT  2.315 2.635 2.545 3.245 ;
      RECT  2.315 3.245 3.53 3.475 ;
      RECT  8.55 0.37 11.93 0.6 ;
      RECT  8.55 0.6 8.78 1.565 ;
      RECT  7.67 1.565 8.78 1.795 ;
      RECT  7.67 1.795 7.9 2.405 ;
      RECT  2.775 2.405 7.9 2.635 ;
      RECT  7.67 2.635 7.9 3.245 ;
      RECT  7.67 3.245 8.78 3.475 ;
      RECT  12.71 0.37 14.17 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  9.97 1.005 12.94 1.235 ;
      RECT  9.97 1.235 10.2 1.565 ;
      RECT  9.035 1.565 10.2 1.795 ;
      RECT  9.035 1.795 9.265 2.405 ;
      RECT  8.23 2.405 9.265 2.635 ;
      RECT  9.035 2.635 9.265 3.245 ;
      RECT  9.035 3.245 10.25 3.475 ;
      RECT  15.27 0.37 18.65 0.6 ;
      RECT  15.27 0.6 15.5 1.565 ;
      RECT  14.39 1.565 15.5 1.795 ;
      RECT  14.39 1.795 14.62 2.405 ;
      RECT  9.495 2.405 14.62 2.635 ;
      RECT  14.39 2.635 14.62 3.245 ;
      RECT  14.39 3.245 15.5 3.475 ;
      RECT  19.385 0.37 20.895 0.6 ;
      RECT  19.385 0.6 19.615 1.005 ;
      RECT  16.7 1.005 19.615 1.235 ;
      RECT  16.7 1.235 16.93 1.565 ;
      RECT  15.755 1.565 16.93 1.795 ;
      RECT  15.755 1.795 15.985 2.405 ;
      RECT  14.905 2.405 15.985 2.635 ;
      RECT  15.755 2.635 15.985 3.245 ;
      RECT  15.755 3.245 16.97 3.475 ;
      RECT  21.99 0.37 25.37 0.6 ;
      RECT  21.99 0.6 22.22 1.565 ;
      RECT  21.11 1.565 22.22 1.795 ;
      RECT  21.11 1.795 21.34 2.38 ;
      RECT  16.215 2.38 21.34 2.61 ;
      RECT  21.11 2.61 21.34 3.245 ;
      RECT  21.11 3.245 22.22 3.475 ;
      RECT  26.105 0.37 27.61 0.6 ;
      RECT  26.105 0.6 26.335 1.005 ;
      RECT  23.405 1.005 26.335 1.235 ;
      RECT  23.405 1.235 23.635 1.565 ;
      RECT  22.475 1.565 23.635 1.795 ;
      RECT  22.475 1.795 22.705 2.405 ;
      RECT  21.67 2.405 22.705 2.635 ;
      RECT  22.475 2.635 22.705 3.245 ;
      RECT  22.475 3.245 23.69 3.475 ;
      RECT  28.71 0.37 32.09 0.6 ;
      RECT  28.71 0.6 28.94 1.565 ;
      RECT  27.83 1.565 28.94 1.795 ;
      RECT  27.83 1.795 28.06 2.41 ;
      RECT  22.935 2.41 28.06 2.64 ;
      RECT  27.83 2.64 28.06 3.245 ;
      RECT  27.83 3.245 28.94 3.475 ;
      RECT  32.865 0.37 34.33 0.6 ;
      RECT  32.865 0.6 33.095 1.005 ;
      RECT  30.125 1.005 33.095 1.235 ;
      RECT  30.125 1.235 30.355 1.565 ;
      RECT  29.195 1.565 30.355 1.795 ;
      RECT  29.195 1.795 29.425 2.405 ;
      RECT  28.39 2.405 29.425 2.635 ;
      RECT  29.195 2.635 29.425 3.245 ;
      RECT  29.195 3.245 30.41 3.475 ;
      RECT  35.43 0.37 38.81 0.6 ;
      RECT  35.43 0.6 35.66 1.565 ;
      RECT  34.55 1.565 35.66 1.795 ;
      RECT  34.55 1.795 34.78 2.405 ;
      RECT  29.655 2.405 34.78 2.635 ;
      RECT  34.55 2.635 34.78 3.245 ;
      RECT  34.55 3.245 35.66 3.475 ;
      RECT  39.59 0.37 41.055 0.6 ;
      RECT  39.59 0.6 39.82 1.005 ;
      RECT  36.9 1.005 39.82 1.235 ;
      RECT  36.9 1.235 37.13 1.565 ;
      RECT  35.915 1.565 37.13 1.795 ;
      RECT  35.915 1.795 36.145 2.405 ;
      RECT  35.065 2.405 36.145 2.635 ;
      RECT  35.915 2.635 36.145 3.245 ;
      RECT  35.915 3.245 37.13 3.475 ;
      RECT  42.15 0.37 45.53 0.6 ;
      RECT  42.15 0.6 42.38 1.565 ;
      RECT  41.27 1.565 42.38 1.795 ;
      RECT  41.27 1.795 41.5 2.375 ;
      RECT  36.385 2.375 41.5 2.605 ;
      RECT  41.27 2.605 41.5 3.245 ;
      RECT  41.27 3.245 42.38 3.475 ;
      RECT  46.3 0.37 47.77 0.6 ;
      RECT  46.3 0.6 46.53 1.005 ;
      RECT  43.565 1.005 46.53 1.235 ;
      RECT  43.565 1.235 43.795 1.565 ;
      RECT  42.7 1.565 43.795 1.795 ;
      RECT  42.7 1.795 42.93 2.405 ;
      RECT  41.825 2.405 42.93 2.635 ;
      RECT  42.7 2.635 42.93 3.245 ;
      RECT  42.7 3.245 43.85 3.475 ;
      RECT  48.87 0.37 52.25 0.6 ;
      RECT  48.87 0.6 49.1 1.565 ;
      RECT  47.99 1.565 49.1 1.795 ;
      RECT  47.99 1.795 48.22 2.41 ;
      RECT  43.16 2.41 48.22 2.64 ;
      RECT  47.99 2.64 48.22 3.245 ;
      RECT  47.99 3.245 49.1 3.475 ;
      RECT  54.13 0.37 54.49 0.6 ;
      RECT  54.13 0.6 54.36 1.005 ;
      RECT  50.34 1.005 54.995 1.235 ;
      RECT  50.34 1.235 50.57 1.565 ;
      RECT  54.765 1.235 54.995 2.405 ;
      RECT  49.44 1.565 50.57 1.795 ;
      RECT  49.44 1.795 49.67 2.405 ;
      RECT  48.55 2.405 49.67 2.635 ;
      RECT  54.765 2.405 55.61 2.635 ;
      RECT  49.44 2.635 49.67 3.245 ;
      RECT  49.44 3.245 50.57 3.475 ;
      RECT  3.95 1.565 5.0 1.795 ;
      RECT  6.185 1.565 7.24 1.795 ;
      RECT  10.67 1.565 11.72 1.795 ;
      RECT  12.92 1.565 13.96 1.795 ;
      RECT  17.39 1.565 18.44 1.795 ;
      RECT  19.625 1.565 20.68 1.795 ;
      RECT  24.11 1.565 25.16 1.795 ;
      RECT  26.345 1.565 27.4 1.795 ;
      RECT  30.84 1.565 31.88 1.795 ;
      RECT  33.065 1.565 34.12 1.795 ;
      RECT  37.56 1.565 38.6 1.795 ;
      RECT  39.8 1.565 40.84 1.795 ;
      RECT  44.27 1.565 45.32 1.795 ;
      RECT  46.505 1.565 47.56 1.795 ;
      RECT  50.99 1.565 52.04 1.795 ;
      RECT  53.835 1.565 54.28 1.795 ;
      RECT  53.835 1.795 54.065 2.405 ;
      RECT  53.17 2.405 54.065 2.635 ;
      RECT  53.835 2.635 54.065 3.245 ;
      RECT  53.835 3.245 54.28 3.475 ;
      RECT  3.96 3.245 5.0 3.475 ;
      RECT  6.165 3.245 7.24 3.475 ;
      RECT  10.68 3.245 11.72 3.475 ;
      RECT  12.92 3.245 13.96 3.475 ;
      RECT  17.4 3.245 18.44 3.475 ;
      RECT  19.605 3.245 20.68 3.475 ;
      RECT  24.12 3.245 25.16 3.475 ;
      RECT  26.325 3.245 27.4 3.475 ;
      RECT  30.84 3.245 31.88 3.475 ;
      RECT  33.045 3.245 34.12 3.475 ;
      RECT  37.56 3.245 38.6 3.475 ;
      RECT  39.8 3.245 40.84 3.475 ;
      RECT  44.28 3.245 45.32 3.475 ;
      RECT  46.485 3.245 47.56 3.475 ;
      RECT  51.0 3.245 52.04 3.475 ;
      RECT  51.95 4.365 53.19 4.37 ;
      RECT  51.95 4.37 53.23 4.595 ;
      RECT  51.95 4.595 52.18 5.0 ;
      RECT  53.0 4.595 53.23 5.0 ;
      RECT  49.67 5.0 52.18 5.23 ;
      RECT  53.0 5.0 53.37 5.23 ;
  END
END MDN_DEL_R64_1
#-----------------------------------------------------------------------
#      Cell        : MDN_DEL_R4_1
#      Description : Delay buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_DEL_R4_1
  CLASS CORE ;
  FOREIGN MDN_DEL_R4_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 1.74 1.235 ;
      RECT  1.005 1.235 1.235 3.245 ;
      RECT  0.18 3.245 1.235 3.475 ;
      RECT  4.11 0.37 5.23 0.6 ;
      RECT  4.11 0.6 4.34 1.565 ;
      RECT  3.96 1.565 4.34 1.795 ;
      RECT  4.11 1.795 4.34 3.245 ;
      RECT  3.96 3.245 4.34 3.475 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  4.715 1.005 6.22 1.235 ;
      RECT  4.715 1.235 4.945 3.5 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.4 ;
      RECT  1.565 2.4 2.76 2.63 ;
      RECT  1.565 2.63 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  2.38 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 2.42 ;
      RECT  3.245 2.42 3.875 2.655 ;
      RECT  3.245 2.655 3.475 3.245 ;
      RECT  2.42 3.245 3.475 3.475 ;
  END
END MDN_DEL_R4_1
#-----------------------------------------------------------------------
#      Cell        : MDN_DEL_R8_1
#      Description : Delay buffer
#      Equation    : X=A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_DEL_R8_1
  CLASS CORE ;
  FOREIGN MDN_DEL_R8_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  6.9 4.365 7.395 4.595 ;
      RECT  7.165 4.595 7.395 5.46 ;
      RECT  6.72 5.46 7.395 5.74 ;
      RECT  4.66 4.365 5.155 4.595 ;
      RECT  4.925 4.595 5.155 5.46 ;
      RECT  4.48 5.46 5.155 5.74 ;
      RECT  2.42 4.365 2.915 4.595 ;
      RECT  2.685 4.595 2.915 5.46 ;
      RECT  2.24 5.46 2.915 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  5.04 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 1.005 ;
      RECT  4.66 1.005 7.255 1.235 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.14 1.005 2.76 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.525 1.565 11.02 1.795 ;
      RECT  10.525 1.795 10.755 3.245 ;
      RECT  10.525 3.245 11.02 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 5.21 0.6 ;
      RECT  3.245 0.6 3.475 1.565 ;
      RECT  3.245 1.565 4.3 1.795 ;
      RECT  3.245 1.795 3.475 3.245 ;
      RECT  3.245 3.245 4.3 3.475 ;
      RECT  5.99 0.37 7.955 0.6 ;
      RECT  7.725 0.6 7.955 1.565 ;
      RECT  7.725 1.565 8.78 1.795 ;
      RECT  8.285 1.795 8.515 2.41 ;
      RECT  8.285 2.41 9.48 2.64 ;
      RECT  8.285 2.64 8.515 3.245 ;
      RECT  7.67 3.245 8.78 3.475 ;
      RECT  10.425 0.37 10.81 0.6 ;
      RECT  10.425 0.6 10.655 1.005 ;
      RECT  8.23 0.37 8.57 0.6 ;
      RECT  8.34 0.6 8.57 1.005 ;
      RECT  8.34 1.005 10.655 1.235 ;
      RECT  9.965 1.235 10.195 3.245 ;
      RECT  9.14 3.245 10.195 3.475 ;
      RECT  0.95 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.405 ;
      RECT  1.565 2.405 2.76 2.635 ;
      RECT  1.565 2.635 1.795 3.245 ;
      RECT  0.95 3.245 2.065 3.475 ;
      RECT  5.38 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 2.405 ;
      RECT  3.75 2.405 7.285 2.635 ;
      RECT  6.045 2.635 6.275 3.245 ;
      RECT  5.43 3.245 6.54 3.475 ;
  END
END MDN_DEL_R8_1
#-----------------------------------------------------------------------
#      Cell        : MDN_EN2_1
#      Description : 2-Input exclusive NOR
#      Equation    : X=!(A1^A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_EN2_1
  CLASS CORE ;
  FOREIGN MDN_EN2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 4.365 5.18 5.0 ;
      RECT  2.63 5.0 5.19 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 1.51 3.475 3.53 ;
    END
    ANTENNADIFFAREA 2.566 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.565 0.445 4.035 0.675 ;
      RECT  1.565 0.675 1.795 1.005 ;
      RECT  3.805 0.675 4.035 1.005 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  1.565 1.565 2.76 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 3.475 4.035 ;
      RECT  3.245 4.035 3.475 4.365 ;
      RECT  3.245 4.365 4.3 4.595 ;
      RECT  4.365 1.565 5.0 1.795 ;
      RECT  4.365 1.795 4.595 2.405 ;
      RECT  3.75 2.405 4.595 2.635 ;
      RECT  4.365 2.635 4.595 3.245 ;
      RECT  4.365 3.245 5.0 3.475 ;
  END
END MDN_EN2_1
#-----------------------------------------------------------------------
#      Cell        : MDN_EN2_2
#      Description : 2-Input exclusive NOR
#      Equation    : X=!(A1^A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_EN2_2
  CLASS CORE ;
  FOREIGN MDN_EN2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  6.2 3.245 7.24 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.19 1.005 6.22 1.235 ;
      RECT  5.485 1.235 5.715 3.805 ;
      RECT  3.19 3.805 5.715 4.035 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  1.565 1.565 4.3 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 2.76 4.035 ;
      RECT  4.715 1.51 4.945 2.405 ;
      RECT  3.75 2.405 4.945 2.635 ;
      RECT  4.715 2.635 4.945 3.53 ;
      RECT  2.63 5.0 5.21 5.23 ;
  END
END MDN_EN2_2
#-----------------------------------------------------------------------
#      Cell        : MDN_EN2_3
#      Description : 2-Input exclusive NOR
#      Equation    : X=!(A1^A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_EN2_3
  CLASS CORE ;
  FOREIGN MDN_EN2_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 8.78 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  6.2 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 4.536 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  3.19 1.005 5.715 1.235 ;
      RECT  5.485 1.235 5.715 2.405 ;
      RECT  5.485 2.405 6.235 2.635 ;
      RECT  5.485 2.635 5.715 3.805 ;
      RECT  3.14 3.805 5.715 4.035 ;
      RECT  1.525 1.565 4.3 1.795 ;
      RECT  1.525 1.795 1.755 3.805 ;
      RECT  1.525 3.805 2.76 4.035 ;
      RECT  4.715 1.655 4.945 2.38 ;
      RECT  3.75 2.38 4.945 2.61 ;
      RECT  4.715 2.61 4.945 3.38 ;
      RECT  7.23 2.43 8.57 2.66 ;
      RECT  2.63 5.0 5.21 5.23 ;
  END
END MDN_EN2_3
#-----------------------------------------------------------------------
#      Cell        : MDN_EN2_4
#      Description : 2-Input exclusive NOR
#      Equation    : X=!(A1^A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_EN2_4
  CLASS CORE ;
  FOREIGN MDN_EN2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 10.195 1.795 ;
      RECT  9.965 1.795 10.195 3.245 ;
      RECT  6.2 3.245 10.195 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  1.505 4.595 1.735 5.0 ;
      RECT  1.505 5.0 1.85 5.23 ;
      RECT  3.19 1.005 5.715 1.235 ;
      RECT  5.485 1.235 5.715 2.405 ;
      RECT  5.485 2.405 9.565 2.635 ;
      RECT  5.485 2.635 5.715 3.805 ;
      RECT  3.19 3.805 5.715 4.035 ;
      RECT  1.565 1.565 4.3 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 2.76 4.035 ;
      RECT  4.66 1.565 5.0 1.795 ;
      RECT  4.66 1.795 4.89 2.375 ;
      RECT  3.75 2.375 4.89 2.605 ;
      RECT  4.66 2.605 4.89 3.245 ;
      RECT  4.66 3.245 5.0 3.475 ;
      RECT  2.63 5.0 5.21 5.23 ;
  END
END MDN_EN2_4
#-----------------------------------------------------------------------
#      Cell        : MDN_EN3_1
#      Description : 3-Input exclusive NOR
#      Equation    : X=!((A1^A2)^A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_EN3_1
  CLASS CORE ;
  FOREIGN MDN_EN3_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.23 0.37 11.34 0.6 ;
      RECT  11.06 0.6 11.34 1.235 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.11 0.37 7.45 0.6 ;
      RECT  7.14 0.6 7.42 1.235 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  7.725 5.02 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  1.005 5.02 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.765 1.565 13.26 1.795 ;
      RECT  12.765 1.795 12.995 3.245 ;
      RECT  12.765 3.245 13.26 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 6.54 1.235 ;
      RECT  2.63 0.37 6.33 0.6 ;
      RECT  9.955 1.005 10.445 1.235 ;
      RECT  10.215 1.235 10.445 3.445 ;
      RECT  9.91 3.445 10.445 3.675 ;
      RECT  4.365 1.565 5.0 1.795 ;
      RECT  4.365 1.795 4.595 3.555 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.555 ;
      RECT  2.685 3.555 6.485 3.785 ;
      RECT  6.255 3.19 6.485 3.555 ;
      RECT  2.685 3.785 2.915 3.805 ;
      RECT  1.72 3.805 2.915 4.035 ;
      RECT  9.14 1.565 9.985 1.795 ;
      RECT  9.755 1.795 9.985 2.965 ;
      RECT  9.26 2.965 9.985 3.195 ;
      RECT  9.26 3.195 9.49 4.015 ;
      RECT  3.24 4.015 10.965 4.245 ;
      RECT  10.735 3.75 10.965 4.015 ;
      RECT  10.675 1.565 11.43 1.795 ;
      RECT  11.2 1.795 11.43 4.475 ;
      RECT  5.43 4.475 11.43 4.705 ;
      RECT  8.495 1.51 8.725 2.36 ;
      RECT  8.495 2.36 9.525 2.59 ;
      RECT  8.495 2.59 8.725 3.53 ;
      RECT  6.955 1.63 7.185 2.405 ;
      RECT  5.99 2.405 7.185 2.635 ;
      RECT  6.955 2.635 7.185 3.53 ;
      RECT  3.245 1.51 3.475 3.315 ;
      RECT  5.485 1.51 5.715 3.315 ;
      RECT  11.72 4.365 12.94 4.595 ;
      RECT  11.72 4.595 11.95 4.985 ;
      RECT  12.71 4.595 12.94 5.0 ;
      RECT  9.91 4.985 11.95 5.215 ;
      RECT  12.71 5.0 13.05 5.23 ;
      RECT  0.18 4.48 5.0 4.71 ;
      RECT  1.51 4.71 1.74 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  3.75 5.0 7.45 5.23 ;
  END
END MDN_EN3_1
#-----------------------------------------------------------------------
#      Cell        : MDN_EN3_2
#      Description : 3-Input exclusive NOR
#      Equation    : X=!((A1^A2)^A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_EN3_2
  CLASS CORE ;
  FOREIGN MDN_EN3_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.23 0.37 9.69 0.6 ;
      RECT  8.26 0.6 8.54 1.235 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  7.725 5.025 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.38 1.565 13.26 1.795 ;
      RECT  12.205 1.795 12.435 2.685 ;
      RECT  11.38 2.685 12.435 2.915 ;
      RECT  12.205 2.915 12.435 3.245 ;
      RECT  11.38 2.915 11.745 3.305 ;
      RECT  12.205 3.245 13.26 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 6.54 1.235 ;
      RECT  3.75 0.37 7.45 0.6 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  11.59 0.37 11.93 0.6 ;
      RECT  11.7 0.6 11.93 1.005 ;
      RECT  9.965 1.005 12.94 1.235 ;
      RECT  9.965 1.235 10.195 3.315 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 3.55 ;
      RECT  1.72 1.565 2.76 1.795 ;
      RECT  2.125 1.795 2.355 3.245 ;
      RECT  1.72 3.245 2.355 3.475 ;
      RECT  2.125 3.475 2.355 3.55 ;
      RECT  2.125 3.55 5.46 3.78 ;
      RECT  5.23 3.78 5.46 4.01 ;
      RECT  5.23 4.01 6.54 4.24 ;
      RECT  10.525 1.565 11.02 1.795 ;
      RECT  10.525 1.795 10.755 3.56 ;
      RECT  10.525 3.56 11.505 3.79 ;
      RECT  11.275 3.79 11.505 4.54 ;
      RECT  7.725 4.005 9.425 4.235 ;
      RECT  7.725 4.235 7.955 4.47 ;
      RECT  9.195 4.235 9.425 4.54 ;
      RECT  3.19 4.47 7.955 4.7 ;
      RECT  9.195 4.54 11.505 4.77 ;
      RECT  6.955 1.54 7.185 2.405 ;
      RECT  5.99 2.405 7.185 2.635 ;
      RECT  6.955 2.635 7.185 3.315 ;
      RECT  5.485 1.51 5.715 3.085 ;
      RECT  5.485 3.085 6.67 3.315 ;
      RECT  6.44 3.315 6.67 3.545 ;
      RECT  6.44 3.545 9.93 3.775 ;
      RECT  9.195 1.585 9.425 3.545 ;
      RECT  9.7 3.775 9.93 4.025 ;
      RECT  9.7 4.025 11.02 4.255 ;
      RECT  3.245 1.51 3.475 3.09 ;
      RECT  3.19 3.09 3.53 3.32 ;
      RECT  8.495 1.54 8.725 3.315 ;
      RECT  1.51 4.01 5.0 4.24 ;
      RECT  1.51 4.24 1.74 4.365 ;
      RECT  0.18 4.365 1.74 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  8.44 4.48 8.78 4.71 ;
      RECT  8.55 4.71 8.78 5.0 ;
      RECT  8.55 5.0 10.81 5.23 ;
      RECT  2.63 5.0 6.33 5.23 ;
  END
END MDN_EN3_2
#-----------------------------------------------------------------------
#      Cell        : MDN_EN3_4
#      Description : 3-Input exclusive NOR
#      Equation    : X=!((A1^A2)^A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_EN3_4
  CLASS CORE ;
  FOREIGN MDN_EN3_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.23 0.37 9.69 0.6 ;
      RECT  8.26 0.6 8.54 1.235 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  7.725 5.02 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.38 1.565 15.5 1.795 ;
      RECT  12.205 1.795 12.435 2.685 ;
      RECT  11.38 2.685 12.435 2.915 ;
      RECT  12.205 2.915 12.435 3.245 ;
      RECT  11.38 2.915 11.72 3.27 ;
      RECT  12.205 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 6.545 1.235 ;
      RECT  3.75 0.37 7.45 0.6 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  11.59 0.37 11.93 0.6 ;
      RECT  11.7 0.6 11.93 1.005 ;
      RECT  9.965 1.005 12.94 1.235 ;
      RECT  9.965 1.235 10.195 3.375 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 3.55 ;
      RECT  1.72 1.565 2.76 1.795 ;
      RECT  2.125 1.795 2.355 3.55 ;
      RECT  1.72 3.55 5.715 3.78 ;
      RECT  5.485 3.78 5.715 4.015 ;
      RECT  5.485 4.015 6.54 4.245 ;
      RECT  6.605 1.565 7.24 1.795 ;
      RECT  6.605 1.795 6.835 2.405 ;
      RECT  5.99 2.405 6.835 2.635 ;
      RECT  6.605 2.635 6.835 3.04 ;
      RECT  6.605 3.04 7.24 3.27 ;
      RECT  10.525 1.565 11.02 1.795 ;
      RECT  10.525 1.795 10.755 3.525 ;
      RECT  10.525 3.525 11.875 3.755 ;
      RECT  11.645 3.755 11.875 4.48 ;
      RECT  7.725 4.02 9.335 4.25 ;
      RECT  7.725 4.25 7.955 4.475 ;
      RECT  9.105 4.25 9.335 4.48 ;
      RECT  3.19 4.475 7.955 4.705 ;
      RECT  9.105 4.48 11.875 4.71 ;
      RECT  12.71 2.405 15.29 2.635 ;
      RECT  5.485 1.505 5.715 3.085 ;
      RECT  5.485 3.085 6.275 3.315 ;
      RECT  6.045 3.315 6.275 3.555 ;
      RECT  6.045 3.555 9.81 3.785 ;
      RECT  9.195 1.58 9.425 3.555 ;
      RECT  9.58 3.785 9.81 4.015 ;
      RECT  9.58 4.015 11.02 4.245 ;
      RECT  3.245 1.51 3.475 3.315 ;
      RECT  8.495 1.585 8.725 3.325 ;
      RECT  1.51 4.01 5.0 4.24 ;
      RECT  1.51 4.24 1.74 4.365 ;
      RECT  0.18 4.365 1.74 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  8.44 4.48 8.78 4.71 ;
      RECT  8.55 4.71 8.78 5.0 ;
      RECT  8.55 5.0 10.81 5.23 ;
      RECT  2.63 5.0 6.33 5.23 ;
  END
END MDN_EN3_4
#-----------------------------------------------------------------------
#      Cell        : MDN_EO2_1
#      Description : 2-Input exclusive OR
#      Equation    : X=A1^A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_EO2_1
  CLASS CORE ;
  FOREIGN MDN_EO2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 4.365 5.18 5.0 ;
      RECT  3.75 5.0 5.21 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.905 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.905 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 1.51 3.475 3.53 ;
    END
    ANTENNADIFFAREA 2.566 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  2.63 0.37 2.97 0.375 ;
      RECT  2.63 0.375 5.155 0.6 ;
      RECT  2.69 0.6 5.155 0.605 ;
      RECT  4.925 0.605 5.155 1.005 ;
      RECT  4.66 1.005 5.155 1.235 ;
      RECT  4.925 1.235 5.155 3.245 ;
      RECT  4.66 3.245 5.155 3.475 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  1.565 1.565 2.76 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 3.475 4.035 ;
      RECT  3.245 4.035 3.475 4.365 ;
      RECT  3.245 4.365 4.3 4.595 ;
  END
END MDN_EO2_1
#-----------------------------------------------------------------------
#      Cell        : MDN_EO2_2
#      Description : 2-Input exclusive OR
#      Equation    : X=A1^A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_EO2_2
  CLASS CORE ;
  FOREIGN MDN_EO2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.195 1.565 7.24 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  6.2 3.245 7.24 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.19 0.445 5.155 0.675 ;
      RECT  4.925 0.675 5.155 1.005 ;
      RECT  4.925 1.005 6.22 1.235 ;
      RECT  5.485 1.235 5.715 4.365 ;
      RECT  3.19 4.365 5.715 4.595 ;
      RECT  1.53 1.565 2.76 1.795 ;
      RECT  1.53 1.795 1.76 3.805 ;
      RECT  1.53 3.805 4.3 4.035 ;
      RECT  4.715 1.585 4.945 2.415 ;
      RECT  3.75 2.415 4.945 2.645 ;
      RECT  4.715 2.645 4.945 3.53 ;
      RECT  2.63 5.0 5.21 5.23 ;
  END
END MDN_EO2_2
#-----------------------------------------------------------------------
#      Cell        : MDN_EO2_3
#      Description : 2-Input exclusive OR
#      Equation    : X=A1^A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_EO2_3
  CLASS CORE ;
  FOREIGN MDN_EO2_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.84 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 8.78 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  6.2 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 4.536 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  3.19 0.445 5.155 0.675 ;
      RECT  4.925 0.675 5.155 1.005 ;
      RECT  4.925 1.005 5.715 1.235 ;
      RECT  5.485 1.235 5.715 2.41 ;
      RECT  5.485 2.41 6.21 2.64 ;
      RECT  5.485 2.64 5.715 4.365 ;
      RECT  3.19 4.365 5.715 4.595 ;
      RECT  1.565 1.565 2.76 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 4.3 4.035 ;
      RECT  4.715 1.585 4.945 2.405 ;
      RECT  3.75 2.405 4.945 2.635 ;
      RECT  4.715 2.635 4.945 3.37 ;
      RECT  7.11 2.405 8.455 2.635 ;
      RECT  2.63 5.0 5.21 5.23 ;
  END
END MDN_EO2_3
#-----------------------------------------------------------------------
#      Cell        : MDN_EO2_4
#      Description : 2-Input exclusive OR
#      Equation    : X=A1^A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_EO2_4
  CLASS CORE ;
  FOREIGN MDN_EO2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 10.195 1.795 ;
      RECT  9.965 1.795 10.195 3.245 ;
      RECT  6.09 3.245 10.195 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  3.19 0.445 5.155 0.675 ;
      RECT  4.925 0.675 5.155 1.005 ;
      RECT  4.925 1.005 5.715 1.235 ;
      RECT  5.485 1.235 5.715 2.405 ;
      RECT  5.485 2.405 9.625 2.635 ;
      RECT  5.485 2.635 5.715 4.365 ;
      RECT  3.19 4.365 5.715 4.595 ;
      RECT  1.53 1.565 2.76 1.795 ;
      RECT  1.53 1.795 1.76 3.805 ;
      RECT  1.53 3.805 4.3 4.035 ;
      RECT  4.715 1.585 4.945 2.415 ;
      RECT  3.75 2.415 4.945 2.645 ;
      RECT  4.715 2.645 4.945 3.37 ;
      RECT  2.63 5.0 5.21 5.23 ;
  END
END MDN_EO2_4
#-----------------------------------------------------------------------
#      Cell        : MDN_EO3_1
#      Description : 3-Input exclusive OR
#      Equation    : X=(A1^A2)^A3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_EO3_1
  CLASS CORE ;
  FOREIGN MDN_EO3_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.23 0.37 9.69 0.6 ;
      RECT  9.38 0.6 9.66 1.235 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.75 0.37 7.45 0.6 ;
      RECT  7.14 0.6 7.42 1.235 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.765 1.565 13.26 1.795 ;
      RECT  12.765 1.795 12.995 3.245 ;
      RECT  12.765 3.245 13.26 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.765 1.48 5.005 1.71 ;
      RECT  3.765 1.71 3.995 3.55 ;
      RECT  1.69 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 3.55 ;
      RECT  1.72 3.55 5.715 3.78 ;
      RECT  5.485 3.545 5.715 3.55 ;
      RECT  5.485 3.78 5.715 4.01 ;
      RECT  5.485 4.01 6.54 4.24 ;
      RECT  10.525 1.565 11.02 1.795 ;
      RECT  10.525 1.795 10.755 2.685 ;
      RECT  10.525 2.685 11.515 2.915 ;
      RECT  11.285 2.915 11.515 4.01 ;
      RECT  7.165 4.01 11.515 4.24 ;
      RECT  7.165 4.24 7.395 4.54 ;
      RECT  3.19 4.54 7.395 4.77 ;
      RECT  5.485 1.505 5.715 1.94 ;
      RECT  4.365 1.94 5.715 2.17 ;
      RECT  4.365 2.17 4.595 3.03 ;
      RECT  4.365 3.03 6.275 3.26 ;
      RECT  6.045 3.26 6.275 3.545 ;
      RECT  6.045 3.545 11.02 3.775 ;
      RECT  9.195 1.585 9.425 3.545 ;
      RECT  6.955 1.645 7.185 2.405 ;
      RECT  4.87 2.405 7.185 2.635 ;
      RECT  6.955 2.635 7.185 3.315 ;
      RECT  3.245 1.51 3.475 3.315 ;
      RECT  8.495 1.585 8.725 3.315 ;
      RECT  9.965 1.54 10.195 3.315 ;
      RECT  2.685 4.01 5.0 4.24 ;
      RECT  2.685 4.24 2.915 4.365 ;
      RECT  0.18 1.005 6.235 1.235 ;
      RECT  6.005 1.235 6.235 1.565 ;
      RECT  1.005 1.235 1.235 2.41 ;
      RECT  6.005 1.565 6.54 1.795 ;
      RECT  1.005 2.41 1.76 2.64 ;
      RECT  1.005 2.64 1.235 4.365 ;
      RECT  0.18 4.365 2.915 4.595 ;
      RECT  11.77 4.11 12.895 4.34 ;
      RECT  11.77 4.34 12.0 4.47 ;
      RECT  12.665 4.34 12.895 5.0 ;
      RECT  9.91 4.47 12.0 4.7 ;
      RECT  12.665 5.0 13.05 5.23 ;
      RECT  8.44 4.48 8.78 4.71 ;
      RECT  8.55 4.71 8.78 5.0 ;
      RECT  8.55 5.0 10.8 5.23 ;
      RECT  2.63 5.0 5.21 5.23 ;
  END
END MDN_EO3_1
#-----------------------------------------------------------------------
#      Cell        : MDN_EO3_2
#      Description : 3-Input exclusive OR
#      Equation    : X=(A1^A2)^A3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_EO3_2
  CLASS CORE ;
  FOREIGN MDN_EO3_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.23 0.37 9.69 0.6 ;
      RECT  8.26 0.6 8.54 1.235 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.6 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.38 1.565 13.26 1.795 ;
      RECT  12.205 1.795 12.435 2.685 ;
      RECT  11.57 2.68 11.875 2.685 ;
      RECT  11.57 2.685 12.995 2.915 ;
      RECT  11.57 2.915 11.875 3.16 ;
      RECT  12.765 2.915 12.995 3.245 ;
      RECT  11.38 3.16 11.875 3.39 ;
      RECT  12.765 3.245 13.26 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.62 0.6 1.85 0.83 ;
      RECT  1.62 0.83 6.38 1.005 ;
      RECT  0.18 1.005 6.38 1.06 ;
      RECT  2.42 1.06 2.76 1.12 ;
      RECT  0.18 1.06 1.85 1.235 ;
      RECT  6.15 1.06 6.38 1.565 ;
      RECT  6.15 1.565 6.54 1.795 ;
      RECT  2.63 0.37 7.185 0.6 ;
      RECT  6.955 0.6 7.185 3.315 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 0.95 ;
      RECT  11.59 0.37 11.93 0.6 ;
      RECT  11.7 0.6 11.93 0.95 ;
      RECT  9.965 0.95 12.94 1.18 ;
      RECT  9.965 1.18 10.195 3.315 ;
      RECT  2.92 1.29 5.155 1.295 ;
      RECT  2.915 1.295 5.155 1.3 ;
      RECT  2.91 1.3 5.155 1.305 ;
      RECT  2.905 1.305 5.155 1.31 ;
      RECT  2.9 1.31 5.155 1.315 ;
      RECT  2.895 1.315 5.155 1.32 ;
      RECT  2.89 1.32 5.155 1.325 ;
      RECT  2.885 1.325 5.155 1.33 ;
      RECT  2.88 1.33 5.155 1.335 ;
      RECT  2.875 1.335 5.155 1.34 ;
      RECT  2.87 1.34 5.155 1.345 ;
      RECT  2.865 1.345 5.155 1.35 ;
      RECT  2.86 1.35 5.155 1.355 ;
      RECT  2.855 1.355 5.155 1.36 ;
      RECT  2.85 1.36 5.155 1.365 ;
      RECT  2.845 1.365 5.155 1.37 ;
      RECT  2.84 1.37 5.155 1.375 ;
      RECT  2.835 1.375 5.155 1.38 ;
      RECT  2.83 1.38 5.155 1.385 ;
      RECT  2.825 1.385 5.155 1.39 ;
      RECT  2.82 1.39 5.155 1.395 ;
      RECT  2.815 1.395 5.155 1.4 ;
      RECT  2.81 1.4 5.155 1.405 ;
      RECT  2.805 1.405 5.155 1.41 ;
      RECT  2.8 1.41 5.155 1.415 ;
      RECT  2.795 1.415 5.155 1.42 ;
      RECT  2.79 1.42 5.155 1.425 ;
      RECT  2.785 1.425 5.155 1.43 ;
      RECT  2.78 1.43 5.155 1.435 ;
      RECT  2.775 1.435 5.155 1.44 ;
      RECT  2.77 1.44 5.155 1.445 ;
      RECT  2.765 1.445 5.155 1.45 ;
      RECT  2.76 1.45 5.155 1.455 ;
      RECT  2.755 1.455 5.155 1.46 ;
      RECT  2.75 1.46 5.155 1.465 ;
      RECT  2.745 1.465 5.155 1.47 ;
      RECT  2.74 1.47 5.155 1.475 ;
      RECT  2.735 1.475 5.155 1.48 ;
      RECT  2.73 1.48 5.155 1.485 ;
      RECT  2.725 1.485 5.155 1.49 ;
      RECT  2.72 1.49 5.155 1.495 ;
      RECT  2.715 1.495 5.155 1.5 ;
      RECT  2.71 1.5 5.155 1.505 ;
      RECT  2.705 1.505 5.155 1.51 ;
      RECT  2.7 1.51 5.155 1.515 ;
      RECT  2.695 1.515 5.155 1.52 ;
      RECT  2.69 1.52 3.055 1.525 ;
      RECT  4.925 1.52 5.155 3.565 ;
      RECT  2.685 1.525 3.05 1.53 ;
      RECT  2.68 1.53 3.045 1.535 ;
      RECT  2.675 1.535 3.04 1.54 ;
      RECT  2.67 1.54 3.035 1.545 ;
      RECT  2.665 1.545 3.03 1.55 ;
      RECT  2.66 1.55 3.025 1.555 ;
      RECT  2.655 1.555 3.02 1.56 ;
      RECT  2.65 1.56 3.015 1.565 ;
      RECT  1.72 1.565 3.01 1.57 ;
      RECT  1.72 1.57 3.005 1.575 ;
      RECT  1.72 1.575 3.0 1.58 ;
      RECT  1.72 1.58 2.995 1.585 ;
      RECT  1.72 1.585 2.99 1.59 ;
      RECT  1.72 1.59 2.985 1.595 ;
      RECT  1.72 1.595 2.98 1.6 ;
      RECT  1.72 1.6 2.975 1.605 ;
      RECT  1.72 1.605 2.97 1.61 ;
      RECT  1.72 1.61 2.965 1.615 ;
      RECT  1.72 1.615 2.96 1.62 ;
      RECT  1.72 1.62 2.955 1.625 ;
      RECT  1.72 1.625 2.95 1.63 ;
      RECT  1.72 1.63 2.945 1.635 ;
      RECT  1.72 1.635 2.94 1.64 ;
      RECT  1.72 1.64 2.935 1.645 ;
      RECT  1.72 1.645 2.93 1.65 ;
      RECT  1.72 1.65 2.925 1.655 ;
      RECT  1.72 1.655 2.92 1.66 ;
      RECT  1.72 1.66 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
      RECT  4.925 3.565 5.715 3.795 ;
      RECT  5.485 3.795 5.715 4.01 ;
      RECT  5.485 4.01 6.54 4.24 ;
      RECT  10.68 1.565 11.02 1.57 ;
      RECT  10.525 1.57 11.02 1.795 ;
      RECT  10.525 1.795 10.755 3.62 ;
      RECT  10.525 3.62 11.505 3.85 ;
      RECT  11.275 3.85 11.505 4.54 ;
      RECT  6.795 4.02 9.425 4.25 ;
      RECT  6.795 4.25 7.025 4.505 ;
      RECT  9.195 4.25 9.425 4.54 ;
      RECT  3.19 4.505 7.025 4.735 ;
      RECT  9.195 4.54 11.505 4.77 ;
      RECT  3.24 1.75 3.58 1.98 ;
      RECT  3.24 1.98 3.47 3.53 ;
      RECT  5.485 1.51 5.715 3.095 ;
      RECT  5.485 3.095 6.275 3.325 ;
      RECT  6.045 3.325 6.275 3.545 ;
      RECT  6.045 3.545 9.905 3.775 ;
      RECT  9.195 1.54 9.425 3.545 ;
      RECT  9.675 3.775 9.905 4.08 ;
      RECT  9.675 4.08 11.02 4.31 ;
      RECT  8.495 1.54 8.725 3.315 ;
      RECT  2.685 4.035 5.0 4.265 ;
      RECT  2.685 4.265 2.915 4.365 ;
      RECT  0.18 4.365 2.915 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  8.44 4.48 8.78 4.71 ;
      RECT  8.55 4.71 8.78 5.0 ;
      RECT  8.55 5.0 10.81 5.23 ;
      RECT  3.75 5.0 7.45 5.23 ;
  END
END MDN_EO3_2
#-----------------------------------------------------------------------
#      Cell        : MDN_EO3_4
#      Description : 3-Input exclusive OR
#      Equation    : X=(A1^A2)^A3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_EO3_4
  CLASS CORE ;
  FOREIGN MDN_EO3_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.23 0.37 9.7 0.6 ;
      RECT  8.26 0.6 8.54 1.235 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  11.76 -0.14 12.435 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.66 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.38 1.565 15.5 1.795 ;
      RECT  12.205 1.795 12.435 2.685 ;
      RECT  11.435 2.685 12.435 2.915 ;
      RECT  12.205 2.915 12.435 3.245 ;
      RECT  11.435 2.915 11.665 3.32 ;
      RECT  12.205 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 0.89 ;
      RECT  0.18 0.89 6.43 1.06 ;
      RECT  2.455 0.83 6.43 0.89 ;
      RECT  0.18 1.06 2.76 1.12 ;
      RECT  6.2 1.06 6.43 1.565 ;
      RECT  6.2 1.565 6.54 1.795 ;
      RECT  2.63 0.37 7.185 0.6 ;
      RECT  6.955 0.6 7.185 3.315 ;
      RECT  14.95 0.37 15.29 0.6 ;
      RECT  14.95 0.6 15.18 1.005 ;
      RECT  13.83 0.37 14.17 0.6 ;
      RECT  13.94 0.6 14.17 1.005 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  11.59 0.37 11.93 0.6 ;
      RECT  11.7 0.6 11.93 1.005 ;
      RECT  9.965 1.005 15.18 1.235 ;
      RECT  9.965 1.235 10.195 3.315 ;
      RECT  3.0 1.29 5.155 1.295 ;
      RECT  2.995 1.295 5.155 1.3 ;
      RECT  2.99 1.3 5.155 1.305 ;
      RECT  2.985 1.305 5.155 1.31 ;
      RECT  2.98 1.31 5.155 1.315 ;
      RECT  2.975 1.315 5.155 1.32 ;
      RECT  2.97 1.32 5.155 1.325 ;
      RECT  2.965 1.325 5.155 1.33 ;
      RECT  2.96 1.33 5.155 1.335 ;
      RECT  2.955 1.335 5.155 1.34 ;
      RECT  2.95 1.34 5.155 1.345 ;
      RECT  2.945 1.345 5.155 1.35 ;
      RECT  1.72 1.35 5.155 1.52 ;
      RECT  1.72 1.52 3.095 1.525 ;
      RECT  4.925 1.52 5.155 3.545 ;
      RECT  1.72 1.525 3.09 1.53 ;
      RECT  1.72 1.53 3.085 1.535 ;
      RECT  1.72 1.535 3.08 1.54 ;
      RECT  1.72 1.54 3.075 1.545 ;
      RECT  1.72 1.545 3.07 1.55 ;
      RECT  1.72 1.55 3.065 1.555 ;
      RECT  1.72 1.555 3.06 1.56 ;
      RECT  1.72 1.56 3.055 1.565 ;
      RECT  1.72 1.565 3.05 1.57 ;
      RECT  1.72 1.57 3.045 1.575 ;
      RECT  1.72 1.575 3.04 1.58 ;
      RECT  2.125 1.58 2.355 3.545 ;
      RECT  1.72 3.545 5.715 3.775 ;
      RECT  5.485 3.775 5.715 4.075 ;
      RECT  5.485 4.075 6.54 4.305 ;
      RECT  10.525 1.565 11.02 1.795 ;
      RECT  10.525 1.795 10.755 3.56 ;
      RECT  10.525 3.56 11.505 3.79 ;
      RECT  11.275 3.79 11.505 4.48 ;
      RECT  6.9 4.02 9.33 4.25 ;
      RECT  9.1 4.25 9.33 4.48 ;
      RECT  6.9 4.25 7.13 4.535 ;
      RECT  9.1 4.48 11.505 4.71 ;
      RECT  3.19 4.535 7.13 4.765 ;
      RECT  3.24 1.75 3.58 1.98 ;
      RECT  3.245 1.98 3.475 3.03 ;
      RECT  3.14 3.03 3.48 3.26 ;
      RECT  5.485 1.51 5.715 3.085 ;
      RECT  5.485 3.085 6.275 3.315 ;
      RECT  6.045 3.315 6.275 3.545 ;
      RECT  6.045 3.545 9.905 3.775 ;
      RECT  9.195 1.585 9.425 3.545 ;
      RECT  9.675 3.775 9.905 4.02 ;
      RECT  9.675 4.02 11.02 4.25 ;
      RECT  8.495 1.585 8.725 3.315 ;
      RECT  2.685 4.015 5.0 4.245 ;
      RECT  2.685 4.245 2.915 4.365 ;
      RECT  0.18 4.365 2.915 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  8.44 4.48 8.78 4.71 ;
      RECT  8.55 4.71 8.78 5.0 ;
      RECT  8.55 5.0 10.81 5.23 ;
      RECT  3.745 5.0 7.45 5.23 ;
  END
END MDN_EO3_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FDN_4
#      Description : D-Flip Flop, neg-edge triggered
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDN_4
  CLASS CORE ;
  FOREIGN MDN_FDN_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 24.64 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 7.42 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  20.34 1.565 24.46 1.795 ;
      RECT  22.285 1.795 22.515 3.245 ;
      RECT  20.34 3.245 24.46 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.86 1.565 19.98 1.795 ;
      RECT  17.805 1.795 18.035 3.245 ;
      RECT  15.86 3.245 19.98 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.81 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 21.84 5.74 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.685 5.46 19.6 5.74 ;
      RECT  18.925 4.87 19.155 5.46 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  4.31 5.46 5.715 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 24.64 5.74 ;
      LAYER VIA12 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  24.23 5.47 24.49 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  18.07 5.47 18.33 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 24.81 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  21.165 0.14 21.395 0.73 ;
      RECT  23.405 0.14 23.635 0.73 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  11.76 -0.14 14.675 0.14 ;
      RECT  12.15 0.14 12.49 0.675 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 24.64 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  20.31 -0.13 20.57 0.13 ;
      RECT  20.87 -0.13 21.13 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  22.55 -0.13 22.81 0.13 ;
      RECT  23.11 -0.13 23.37 0.13 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 5.155 0.6 ;
      RECT  4.925 0.6 5.155 1.005 ;
      RECT  4.925 1.005 7.955 1.235 ;
      RECT  7.725 1.235 7.955 2.44 ;
      RECT  7.725 2.44 8.57 2.67 ;
      RECT  7.725 2.67 7.955 3.245 ;
      RECT  6.9 3.245 7.955 3.475 ;
      RECT  8.23 0.37 10.81 0.6 ;
      RECT  23.91 0.37 24.25 0.6 ;
      RECT  23.91 0.6 24.14 1.005 ;
      RECT  21.67 0.37 23.13 0.6 ;
      RECT  21.67 0.6 21.9 1.005 ;
      RECT  22.9 0.6 23.13 1.005 ;
      RECT  19.445 0.37 20.92 0.6 ;
      RECT  19.445 0.6 19.675 1.005 ;
      RECT  20.69 0.6 20.92 1.005 ;
      RECT  14.95 0.37 15.29 0.6 ;
      RECT  14.95 0.6 15.18 1.005 ;
      RECT  14.445 1.005 19.675 1.235 ;
      RECT  20.69 1.005 21.9 1.235 ;
      RECT  22.9 1.005 24.14 1.235 ;
      RECT  14.445 1.235 14.675 2.125 ;
      RECT  13.885 2.125 14.675 2.355 ;
      RECT  13.885 2.355 14.115 2.765 ;
      RECT  11.38 1.565 12.995 1.795 ;
      RECT  12.765 1.795 12.995 2.765 ;
      RECT  12.765 2.765 14.115 2.995 ;
      RECT  12.765 2.995 12.995 3.245 ;
      RECT  11.38 3.245 12.995 3.475 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  9.14 1.005 13.96 1.235 ;
      RECT  3.96 1.48 5.0 1.71 ;
      RECT  8.44 1.565 9.075 1.795 ;
      RECT  8.845 1.795 9.075 2.41 ;
      RECT  8.845 2.41 9.56 2.64 ;
      RECT  10.525 1.565 11.02 1.795 ;
      RECT  10.525 1.795 10.755 3.805 ;
      RECT  6.195 1.505 6.54 1.735 ;
      RECT  6.31 1.735 6.54 3.245 ;
      RECT  4.87 2.405 5.605 2.635 ;
      RECT  5.375 2.635 5.605 3.245 ;
      RECT  5.375 3.245 6.54 3.475 ;
      RECT  6.31 3.475 6.54 3.805 ;
      RECT  6.31 3.805 10.755 4.035 ;
      RECT  3.245 1.51 3.475 1.94 ;
      RECT  3.245 1.94 6.07 2.17 ;
      RECT  5.84 2.17 6.07 2.685 ;
      RECT  3.245 2.17 3.475 3.53 ;
      RECT  9.965 1.65 10.195 3.53 ;
      RECT  2.42 3.805 5.0 4.035 ;
      RECT  11.085 3.805 13.96 4.035 ;
      RECT  11.085 4.035 11.315 4.365 ;
      RECT  10.68 4.365 11.315 4.595 ;
      RECT  1.72 4.365 4.3 4.595 ;
      RECT  4.925 4.365 9.075 4.595 ;
      RECT  4.925 4.595 5.155 5.0 ;
      RECT  8.845 4.595 9.075 5.0 ;
      RECT  2.63 5.0 5.155 5.23 ;
      RECT  8.845 5.0 9.67 5.23 ;
      RECT  18.42 4.365 19.66 4.595 ;
      RECT  18.42 4.595 18.65 5.0 ;
      RECT  19.43 4.595 19.66 5.0 ;
      RECT  15.005 1.56 15.495 1.565 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 4.365 ;
      RECT  15.005 4.365 17.42 4.595 ;
      RECT  16.18 4.595 16.41 5.0 ;
      RECT  17.19 4.595 17.42 5.0 ;
      RECT  16.07 5.0 16.41 5.23 ;
      RECT  17.19 5.0 18.65 5.23 ;
      RECT  19.43 5.0 19.77 5.23 ;
      RECT  9.91 4.925 11.93 5.155 ;
      RECT  11.59 5.155 11.93 5.23 ;
  END
END MDN_FDN_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FDN_1
#      Description : D-Flip Flop, neg-edge triggered
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDN_1
  CLASS CORE ;
  FOREIGN MDN_FDN_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 7.42 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 3.245 ;
      RECT  15.005 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.62 1.565 14.115 1.795 ;
      RECT  13.885 1.795 14.115 3.245 ;
      RECT  13.62 3.245 14.115 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.93 12.435 5.46 ;
      RECT  12.205 5.46 15.85 5.74 ;
      RECT  14.445 4.93 14.675 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 15.85 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 10.81 0.6 ;
      RECT  8.23 0.6 8.46 1.005 ;
      RECT  3.75 0.37 5.155 0.6 ;
      RECT  4.925 0.6 5.155 1.005 ;
      RECT  4.925 1.005 8.46 1.235 ;
      RECT  7.725 1.235 7.955 2.125 ;
      RECT  7.725 2.125 8.515 2.355 ;
      RECT  8.285 2.355 8.515 3.245 ;
      RECT  6.9 3.245 8.515 3.475 ;
      RECT  14.95 0.37 15.29 0.6 ;
      RECT  14.95 0.6 15.18 1.005 ;
      RECT  12.71 0.37 14.115 0.6 ;
      RECT  13.885 0.6 14.115 1.005 ;
      RECT  13.885 1.005 15.18 1.235 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  9.14 1.005 13.26 1.235 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  8.44 1.565 9.635 1.795 ;
      RECT  9.405 1.795 9.635 2.69 ;
      RECT  10.525 1.565 11.02 1.795 ;
      RECT  10.525 1.795 10.755 3.805 ;
      RECT  5.325 1.565 6.63 1.795 ;
      RECT  5.325 1.795 5.555 2.405 ;
      RECT  6.4 1.795 6.63 3.805 ;
      RECT  4.87 2.405 5.555 2.635 ;
      RECT  6.2 3.805 10.755 4.035 ;
      RECT  11.38 1.565 11.875 1.795 ;
      RECT  11.645 1.795 11.875 2.405 ;
      RECT  11.645 2.405 13.05 2.635 ;
      RECT  11.645 2.635 11.875 3.245 ;
      RECT  11.38 3.245 11.875 3.475 ;
      RECT  3.245 1.54 3.475 3.245 ;
      RECT  3.245 3.245 6.05 3.475 ;
      RECT  5.82 2.35 6.05 3.245 ;
      RECT  9.965 1.51 10.195 3.53 ;
      RECT  2.42 3.805 5.0 4.035 ;
      RECT  11.085 3.805 13.26 4.035 ;
      RECT  11.085 4.035 11.315 4.365 ;
      RECT  10.68 4.365 11.315 4.595 ;
      RECT  1.72 4.365 4.3 4.595 ;
      RECT  4.925 4.365 9.075 4.595 ;
      RECT  4.925 4.595 5.155 5.0 ;
      RECT  8.845 4.595 9.075 5.0 ;
      RECT  2.63 5.0 5.155 5.23 ;
      RECT  8.845 5.0 9.69 5.23 ;
      RECT  11.725 4.365 12.995 4.595 ;
      RECT  11.725 4.595 11.955 5.0 ;
      RECT  12.765 4.595 12.995 5.0 ;
      RECT  9.965 4.31 10.195 5.0 ;
      RECT  9.965 5.0 11.955 5.23 ;
      RECT  12.765 5.0 14.17 5.23 ;
  END
END MDN_FDN_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FDN_2
#      Description : D-Flip Flop, neg-edge triggered
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDN_2
  CLASS CORE ;
  FOREIGN MDN_FDN_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 7.42 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.61 1.565 15.5 1.795 ;
      RECT  14.445 1.795 14.675 3.245 ;
      RECT  13.62 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.86 1.565 17.75 1.795 ;
      RECT  16.685 1.795 16.915 3.245 ;
      RECT  15.86 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  12.205 5.46 18.09 5.74 ;
      RECT  14.445 4.87 14.675 5.46 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  12.205 -0.14 15.12 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 10.81 0.6 ;
      RECT  8.23 0.6 8.46 1.005 ;
      RECT  3.75 0.37 5.155 0.6 ;
      RECT  4.925 0.6 5.155 1.005 ;
      RECT  4.925 1.005 8.46 1.235 ;
      RECT  7.725 1.235 7.955 2.12 ;
      RECT  7.725 2.12 8.475 2.35 ;
      RECT  8.245 2.35 8.475 3.24 ;
      RECT  6.91 3.24 8.475 3.245 ;
      RECT  6.9 3.245 8.475 3.47 ;
      RECT  6.9 3.47 7.24 3.475 ;
      RECT  14.95 0.37 15.29 0.6 ;
      RECT  14.95 0.6 15.18 1.005 ;
      RECT  12.71 0.37 14.17 0.6 ;
      RECT  13.94 0.6 14.17 1.005 ;
      RECT  13.94 1.005 15.18 1.235 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  9.14 1.005 13.26 1.235 ;
      RECT  3.96 1.465 5.0 1.695 ;
      RECT  8.44 1.565 9.635 1.795 ;
      RECT  9.405 1.795 9.635 2.69 ;
      RECT  10.485 1.565 11.02 1.795 ;
      RECT  10.485 1.795 10.715 3.805 ;
      RECT  6.2 1.47 6.545 1.7 ;
      RECT  6.315 1.7 6.545 3.245 ;
      RECT  4.87 2.395 5.59 2.625 ;
      RECT  5.36 2.625 5.59 3.245 ;
      RECT  5.36 3.245 6.545 3.475 ;
      RECT  6.315 3.475 6.545 3.805 ;
      RECT  6.315 3.805 10.715 4.035 ;
      RECT  11.38 1.565 11.86 1.795 ;
      RECT  11.63 1.795 11.86 2.685 ;
      RECT  11.63 2.685 12.995 2.915 ;
      RECT  12.765 2.35 12.995 2.685 ;
      RECT  11.63 2.915 11.86 3.245 ;
      RECT  11.38 3.245 11.86 3.475 ;
      RECT  3.245 1.51 3.475 1.93 ;
      RECT  3.245 1.93 6.085 2.16 ;
      RECT  5.855 2.16 6.085 2.685 ;
      RECT  3.245 2.16 3.475 3.53 ;
      RECT  9.965 1.51 10.195 3.53 ;
      RECT  2.42 3.805 5.0 4.035 ;
      RECT  11.04 3.805 13.26 4.035 ;
      RECT  11.04 4.035 11.31 4.365 ;
      RECT  10.68 4.365 11.31 4.595 ;
      RECT  1.715 4.365 4.3 4.595 ;
      RECT  4.925 4.365 9.075 4.595 ;
      RECT  4.925 4.595 5.155 5.0 ;
      RECT  8.845 4.595 9.075 5.0 ;
      RECT  2.63 5.0 5.155 5.23 ;
      RECT  8.845 5.0 9.69 5.23 ;
      RECT  16.175 4.365 17.42 4.595 ;
      RECT  16.175 4.595 16.405 4.925 ;
      RECT  17.19 4.595 17.42 5.0 ;
      RECT  11.7 4.365 15.235 4.595 ;
      RECT  15.005 4.595 15.235 4.925 ;
      RECT  11.7 4.595 11.93 5.0 ;
      RECT  15.005 4.925 16.405 5.0 ;
      RECT  9.965 4.385 10.195 5.0 ;
      RECT  9.965 5.0 11.93 5.23 ;
      RECT  15.005 5.0 16.41 5.155 ;
      RECT  17.19 5.0 17.53 5.23 ;
      RECT  16.07 5.155 16.41 5.23 ;
  END
END MDN_FDN_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNQ_1
#      Description : D-Flip Flop, neg-edge triggered
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNQ_1
  CLASS CORE ;
  FOREIGN MDN_FDNQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.765 1.565 13.26 1.795 ;
      RECT  12.765 1.795 12.995 3.245 ;
      RECT  12.765 3.245 13.26 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 3.475 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.52 ;
      RECT  -0.17 -0.14 3.92 0.14 ;
      RECT  3.19 0.14 3.53 0.465 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  8.845 0.37 10.81 0.6 ;
      RECT  8.845 0.6 9.075 0.75 ;
      RECT  3.805 0.37 7.395 0.6 ;
      RECT  3.805 0.6 4.035 0.695 ;
      RECT  7.165 0.6 7.395 0.75 ;
      RECT  1.565 0.695 4.035 0.925 ;
      RECT  7.165 0.75 9.075 0.98 ;
      RECT  1.565 0.925 2.06 1.125 ;
      RECT  1.565 1.125 1.795 3.805 ;
      RECT  1.565 3.805 2.06 4.035 ;
      RECT  11.085 0.37 11.94 0.6 ;
      RECT  11.085 0.6 11.315 1.005 ;
      RECT  9.91 1.005 11.315 1.235 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  11.645 1.005 12.94 1.235 ;
      RECT  11.645 1.235 11.875 1.565 ;
      RECT  11.38 1.565 11.875 1.795 ;
      RECT  11.645 1.795 11.875 2.405 ;
      RECT  8.23 2.405 11.875 2.635 ;
      RECT  11.645 2.635 11.875 3.245 ;
      RECT  11.38 3.245 11.875 3.475 ;
      RECT  4.365 1.005 6.54 1.18 ;
      RECT  2.42 1.18 6.54 1.235 ;
      RECT  2.42 1.235 4.595 1.41 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 9.075 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  4.97 4.595 5.2 5.0 ;
      RECT  8.845 4.595 9.075 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  4.86 5.0 5.2 5.23 ;
      RECT  8.845 5.0 9.68 5.23 ;
      RECT  6.9 1.21 9.48 1.44 ;
      RECT  7.725 1.44 7.955 3.245 ;
      RECT  3.92 2.405 6.275 2.635 ;
      RECT  6.045 2.635 6.275 3.245 ;
      RECT  6.045 3.245 11.02 3.475 ;
      RECT  5.43 1.565 6.24 1.795 ;
      RECT  6.01 1.795 6.24 1.845 ;
      RECT  6.01 1.845 7.395 2.075 ;
      RECT  7.165 2.075 7.395 2.69 ;
      RECT  3.96 1.64 5.0 1.87 ;
      RECT  8.44 1.75 11.025 1.98 ;
      RECT  3.96 3.245 5.715 3.475 ;
      RECT  5.485 3.475 5.715 3.805 ;
      RECT  5.485 3.805 6.54 4.035 ;
      RECT  2.42 3.805 5.0 4.035 ;
      RECT  8.435 3.805 9.495 4.035 ;
      RECT  5.43 5.0 7.45 5.23 ;
      RECT  9.91 5.0 11.935 5.23 ;
  END
END MDN_FDNQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNQ_2
#      Description : D-Flip Flop, neg-edge triggered
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNQ_2
  CLASS CORE ;
  FOREIGN MDN_FDNQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.765 1.565 13.965 1.795 ;
      RECT  12.765 1.795 12.995 3.245 ;
      RECT  12.765 3.245 13.96 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.03 5.46 12.435 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.52 ;
      RECT  -0.17 -0.14 3.92 0.14 ;
      RECT  3.19 0.14 3.53 0.465 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 10.81 0.445 ;
      RECT  8.845 0.445 10.81 0.675 ;
      RECT  8.845 0.675 9.075 0.75 ;
      RECT  3.805 0.37 7.395 0.6 ;
      RECT  3.805 0.6 4.035 0.695 ;
      RECT  7.165 0.6 7.395 0.75 ;
      RECT  1.775 0.695 4.035 0.925 ;
      RECT  7.165 0.75 9.075 0.98 ;
      RECT  1.775 0.925 2.005 3.53 ;
      RECT  11.085 0.37 11.93 0.6 ;
      RECT  11.085 0.6 11.315 1.005 ;
      RECT  9.91 1.005 11.315 1.235 ;
      RECT  12.71 0.37 14.17 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  11.645 1.005 12.94 1.235 ;
      RECT  11.645 1.235 11.875 1.565 ;
      RECT  11.38 1.565 11.875 1.795 ;
      RECT  11.645 1.795 11.875 2.405 ;
      RECT  8.23 2.405 11.875 2.635 ;
      RECT  11.645 2.635 11.875 3.245 ;
      RECT  11.38 3.245 11.875 3.475 ;
      RECT  4.365 1.005 6.54 1.18 ;
      RECT  2.42 1.18 6.54 1.235 ;
      RECT  2.42 1.235 4.595 1.41 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 9.075 4.595 ;
      RECT  4.97 4.36 5.2 4.365 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  4.97 4.595 5.2 5.0 ;
      RECT  8.845 4.595 9.075 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  4.86 5.0 5.2 5.23 ;
      RECT  8.845 5.0 9.68 5.23 ;
      RECT  6.9 1.21 9.48 1.44 ;
      RECT  7.725 1.44 7.955 3.245 ;
      RECT  3.805 2.155 6.275 2.385 ;
      RECT  3.805 2.385 4.035 2.69 ;
      RECT  6.045 2.385 6.275 3.245 ;
      RECT  6.045 3.245 11.02 3.475 ;
      RECT  3.96 1.64 5.0 1.87 ;
      RECT  5.43 1.695 7.395 1.925 ;
      RECT  7.165 1.925 7.395 2.69 ;
      RECT  8.44 1.745 11.02 1.975 ;
      RECT  4.785 2.615 5.715 2.845 ;
      RECT  4.785 2.845 5.015 3.245 ;
      RECT  5.485 2.845 5.715 3.805 ;
      RECT  3.96 3.245 5.015 3.475 ;
      RECT  5.485 3.805 6.54 4.035 ;
      RECT  2.42 3.805 5.0 4.035 ;
      RECT  8.44 3.805 9.48 4.035 ;
      RECT  5.43 5.0 7.45 5.23 ;
      RECT  9.91 5.0 11.93 5.23 ;
  END
END MDN_FDNQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNQ_4
#      Description : D-Flip Flop, neg-edge triggered
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNQ_4
  CLASS CORE ;
  FOREIGN MDN_FDNQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.765 1.565 16.245 1.795 ;
      RECT  12.765 1.795 12.995 3.245 ;
      RECT  12.765 3.245 16.245 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.03 5.46 12.435 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 3.475 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.205 0.14 12.435 0.735 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.52 ;
      RECT  -0.17 -0.14 3.92 0.14 ;
      RECT  3.19 0.14 3.53 0.545 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  8.845 0.37 10.81 0.6 ;
      RECT  8.845 0.6 9.075 0.75 ;
      RECT  3.805 0.37 7.395 0.6 ;
      RECT  7.165 0.6 7.395 0.75 ;
      RECT  3.805 0.6 4.035 0.83 ;
      RECT  7.165 0.75 9.075 0.98 ;
      RECT  1.565 0.83 4.035 1.06 ;
      RECT  1.565 1.06 2.06 1.235 ;
      RECT  1.565 1.235 1.795 3.805 ;
      RECT  1.565 3.805 2.06 4.035 ;
      RECT  11.085 0.37 11.94 0.6 ;
      RECT  11.085 0.6 11.315 1.005 ;
      RECT  9.91 1.005 11.315 1.235 ;
      RECT  14.95 0.37 16.41 0.6 ;
      RECT  14.95 0.6 15.18 1.005 ;
      RECT  12.71 0.37 14.17 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  13.94 0.6 14.17 1.005 ;
      RECT  11.645 1.005 12.94 1.235 ;
      RECT  13.94 1.005 15.18 1.235 ;
      RECT  11.645 1.235 11.875 1.565 ;
      RECT  11.38 1.565 11.875 1.795 ;
      RECT  11.645 1.795 11.875 2.405 ;
      RECT  8.23 2.405 11.875 2.635 ;
      RECT  11.645 2.635 11.875 3.245 ;
      RECT  11.38 3.245 11.875 3.475 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 9.075 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  4.96 4.595 5.19 5.0 ;
      RECT  8.845 4.595 9.075 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  4.85 5.0 5.19 5.23 ;
      RECT  8.845 5.0 9.69 5.23 ;
      RECT  4.365 1.005 6.54 1.235 ;
      RECT  4.365 1.235 4.595 1.29 ;
      RECT  2.42 1.29 4.595 1.52 ;
      RECT  6.9 1.21 9.48 1.44 ;
      RECT  7.725 1.44 7.955 3.245 ;
      RECT  3.945 2.35 4.175 2.685 ;
      RECT  3.945 2.685 6.265 2.915 ;
      RECT  6.035 2.915 6.265 3.245 ;
      RECT  6.035 3.245 11.02 3.475 ;
      RECT  5.43 1.565 6.275 1.795 ;
      RECT  6.045 1.795 6.275 1.84 ;
      RECT  6.045 1.84 7.395 2.07 ;
      RECT  7.165 2.07 7.395 2.69 ;
      RECT  3.96 1.75 5.0 1.98 ;
      RECT  8.44 1.75 11.02 1.98 ;
      RECT  3.96 3.245 5.715 3.475 ;
      RECT  5.485 3.475 5.715 3.805 ;
      RECT  5.485 3.805 6.54 4.035 ;
      RECT  2.42 3.805 5.0 4.035 ;
      RECT  8.435 3.805 9.495 4.035 ;
      RECT  9.965 4.87 10.195 5.0 ;
      RECT  9.965 5.0 11.93 5.23 ;
      RECT  5.43 5.0 7.45 5.23 ;
  END
END MDN_FDNQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNRB_4
#      Description : D-Flip Flop, neg-edge triggered, lo-async-clear
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNRB_4
  CLASS CORE ;
  FOREIGN MDN_FDNRB_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 24.64 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.095 0.7 2.885 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.15 1.565 18.44 1.795 ;
      RECT  17.805 1.795 18.035 3.245 ;
      RECT  15.16 3.245 18.44 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  20.34 1.565 24.46 1.795 ;
      RECT  22.285 1.795 22.515 3.245 ;
      RECT  20.34 3.245 24.46 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END QN
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.33 1.565 9.66 1.93 ;
      RECT  7.165 1.93 9.66 2.16 ;
      RECT  9.38 2.16 9.66 2.62 ;
      RECT  7.165 2.16 7.395 2.63 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.81 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 21.84 5.74 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.685 5.46 19.155 5.74 ;
      RECT  18.925 4.87 19.155 5.46 ;
      RECT  14.445 4.91 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  9.405 4.925 10.25 5.155 ;
      RECT  9.405 5.155 9.635 5.46 ;
      RECT  7.67 4.925 8.515 5.155 ;
      RECT  8.285 5.155 8.515 5.46 ;
      RECT  8.285 5.46 9.635 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 3.475 5.74 ;
      RECT  3.245 4.92 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 24.64 5.74 ;
      LAYER VIA12 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  24.23 5.47 24.49 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  18.07 5.47 18.33 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 -0.14 24.81 0.14 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  18.925 -0.14 21.395 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  8.79 -0.14 9.52 0.14 ;
      RECT  8.845 0.14 9.075 0.93 ;
      RECT  8.845 0.93 9.48 1.16 ;
      RECT  6.16 -0.14 6.89 0.14 ;
      RECT  6.605 0.14 6.835 0.89 ;
      RECT  6.605 0.89 7.24 1.12 ;
      RECT  -0.17 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.52 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 24.64 0.14 ;
      LAYER VIA12 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  20.31 -0.13 20.57 0.13 ;
      RECT  20.87 -0.13 21.13 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 2.915 0.6 ;
      RECT  2.685 0.6 2.915 0.83 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  2.685 0.83 6.35 1.06 ;
      RECT  6.0 0.37 6.35 0.83 ;
      RECT  0.18 1.005 1.74 1.235 ;
      RECT  5.97 1.06 6.35 1.26 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 1.235 4.595 ;
      RECT  3.75 0.37 5.77 0.6 ;
      RECT  9.965 0.37 13.05 0.6 ;
      RECT  9.965 0.6 10.195 0.98 ;
      RECT  9.89 0.98 10.27 1.26 ;
      RECT  21.67 0.37 23.13 0.6 ;
      RECT  11.38 1.005 13.96 1.235 ;
      RECT  2.42 1.29 5.0 1.52 ;
      RECT  6.605 1.47 8.78 1.565 ;
      RECT  6.2 1.565 8.78 1.7 ;
      RECT  6.2 1.7 6.835 1.795 ;
      RECT  19.485 1.56 19.98 1.79 ;
      RECT  19.485 1.79 19.715 2.385 ;
      RECT  19.485 2.385 21.98 2.615 ;
      RECT  19.485 2.615 19.715 3.245 ;
      RECT  19.485 3.245 19.98 3.475 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 4.46 ;
      RECT  1.565 4.46 11.82 4.69 ;
      RECT  4.98 4.69 5.21 5.0 ;
      RECT  11.59 4.69 11.82 5.0 ;
      RECT  4.87 5.0 5.21 5.23 ;
      RECT  11.59 5.0 11.93 5.23 ;
      RECT  9.965 1.565 11.02 1.795 ;
      RECT  9.965 1.795 10.195 3.07 ;
      RECT  9.14 3.07 10.195 3.3 ;
      RECT  12.765 1.565 13.26 1.795 ;
      RECT  12.765 1.795 12.995 3.53 ;
      RECT  3.245 1.75 5.155 1.98 ;
      RECT  4.925 1.98 5.155 2.125 ;
      RECT  3.245 1.98 3.475 3.49 ;
      RECT  4.925 2.125 6.275 2.355 ;
      RECT  6.045 2.355 6.275 2.86 ;
      RECT  6.045 2.86 8.515 3.09 ;
      RECT  8.285 2.39 8.515 2.86 ;
      RECT  8.285 3.09 8.515 3.53 ;
      RECT  3.245 3.49 4.3 3.72 ;
      RECT  8.28 3.53 12.995 3.76 ;
      RECT  22.82 2.37 24.25 2.6 ;
      RECT  3.805 2.355 4.035 3.03 ;
      RECT  3.805 3.03 5.77 3.26 ;
      RECT  10.525 2.385 10.755 3.03 ;
      RECT  10.525 3.03 12.49 3.26 ;
      RECT  12.205 1.51 12.435 3.03 ;
      RECT  4.66 3.49 7.13 3.72 ;
      RECT  6.9 3.72 7.13 3.99 ;
      RECT  6.9 3.99 8.78 4.22 ;
      RECT  2.42 3.95 6.54 4.18 ;
      RECT  12.92 3.99 13.965 4.22 ;
      RECT  18.42 4.365 19.66 4.595 ;
      RECT  18.42 4.595 18.65 5.0 ;
      RECT  19.43 4.595 19.66 5.0 ;
      RECT  16.2 4.385 17.42 4.615 ;
      RECT  16.2 4.615 16.43 5.0 ;
      RECT  17.19 4.615 17.42 5.0 ;
      RECT  9.14 4.0 12.435 4.23 ;
      RECT  12.205 4.23 12.435 4.45 ;
      RECT  12.205 4.45 15.18 4.68 ;
      RECT  13.94 4.68 14.17 5.0 ;
      RECT  14.95 4.68 15.18 5.0 ;
      RECT  13.83 5.0 14.17 5.23 ;
      RECT  14.95 5.0 16.43 5.23 ;
      RECT  17.19 5.0 18.65 5.23 ;
      RECT  19.43 5.0 19.77 5.23 ;
      LAYER METAL2 ;
      RECT  5.97 0.98 10.27 1.26 ;
      LAYER VIA12 ;
      RECT  6.03 0.99 6.29 1.25 ;
      RECT  9.95 0.99 10.21 1.25 ;
  END
END MDN_FDNRB_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNRB_1
#      Description : D-Flip Flop, neg-edge triggered, lo-async-clear
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNRB_1
  CLASS CORE ;
  FOREIGN MDN_FDNRB_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.86 1.565 16.915 1.795 ;
      RECT  16.685 1.795 16.915 3.245 ;
      RECT  15.86 3.245 16.915 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.245 1.565 17.74 1.795 ;
      RECT  17.245 1.795 17.475 3.245 ;
      RECT  17.245 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END QN
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.885 2.35 14.115 3.245 ;
      RECT  12.205 3.245 14.115 3.475 ;
      RECT  13.885 3.475 14.115 3.48 ;
      RECT  12.205 3.475 12.435 4.02 ;
      RECT  7.17 2.405 7.955 2.635 ;
      RECT  7.725 2.635 7.955 3.755 ;
      RECT  2.66 2.125 2.94 3.755 ;
      RECT  2.66 3.755 9.24 3.985 ;
      RECT  9.01 3.985 9.24 4.02 ;
      RECT  9.01 4.02 12.435 4.25 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.895 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.895 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  12.205 4.94 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  7.67 5.135 8.01 5.46 ;
      RECT  7.28 5.46 8.4 5.74 ;
      RECT  3.19 5.135 3.53 5.46 ;
      RECT  2.8 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.58 ;
      RECT  12.205 -0.14 14.115 0.14 ;
      RECT  12.205 0.14 12.435 0.6 ;
      RECT  13.885 0.14 14.115 0.89 ;
      RECT  13.62 0.89 14.115 1.12 ;
      RECT  6.55 -0.14 7.28 0.14 ;
      RECT  7.01 0.14 7.24 0.89 ;
      RECT  6.9 0.89 7.24 1.12 ;
      RECT  2.07 -0.14 2.915 0.14 ;
      RECT  2.685 0.14 2.915 1.005 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 1.74 1.235 ;
      RECT  3.22 0.37 6.33 0.6 ;
      RECT  3.22 0.6 3.45 1.565 ;
      RECT  1.565 1.565 3.45 1.795 ;
      RECT  1.565 1.795 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  9.01 0.37 11.93 0.6 ;
      RECT  9.01 0.6 9.24 1.225 ;
      RECT  9.005 1.225 9.24 1.23 ;
      RECT  9.0 1.23 9.24 1.235 ;
      RECT  8.995 1.235 9.24 1.24 ;
      RECT  8.99 1.24 9.24 1.245 ;
      RECT  8.985 1.245 9.24 1.25 ;
      RECT  8.98 1.25 9.24 1.255 ;
      RECT  8.975 1.255 9.24 1.26 ;
      RECT  8.97 1.26 9.24 1.265 ;
      RECT  8.965 1.265 9.24 1.27 ;
      RECT  8.96 1.27 9.24 1.275 ;
      RECT  8.955 1.275 9.24 1.28 ;
      RECT  8.95 1.28 9.24 1.285 ;
      RECT  8.945 1.285 9.24 1.29 ;
      RECT  8.94 1.29 9.24 1.295 ;
      RECT  8.935 1.295 9.24 1.3 ;
      RECT  8.93 1.3 9.24 1.305 ;
      RECT  8.925 1.305 9.24 1.31 ;
      RECT  8.92 1.31 9.24 1.315 ;
      RECT  8.915 1.315 9.24 1.32 ;
      RECT  8.91 1.32 9.235 1.325 ;
      RECT  8.905 1.325 9.23 1.33 ;
      RECT  8.9 1.33 9.225 1.335 ;
      RECT  8.895 1.335 9.22 1.34 ;
      RECT  8.89 1.34 9.215 1.345 ;
      RECT  8.885 1.345 9.21 1.35 ;
      RECT  8.285 1.35 9.205 1.355 ;
      RECT  8.285 1.355 9.2 1.36 ;
      RECT  8.285 1.36 9.195 1.365 ;
      RECT  8.285 1.365 9.19 1.37 ;
      RECT  8.285 1.37 9.185 1.375 ;
      RECT  8.285 1.375 9.18 1.38 ;
      RECT  8.285 1.38 9.175 1.385 ;
      RECT  8.285 1.385 9.17 1.39 ;
      RECT  8.285 1.39 9.165 1.395 ;
      RECT  8.285 1.395 9.16 1.4 ;
      RECT  8.285 1.4 9.155 1.405 ;
      RECT  8.285 1.405 9.15 1.41 ;
      RECT  8.285 1.41 9.145 1.415 ;
      RECT  8.285 1.415 9.14 1.42 ;
      RECT  8.285 1.42 9.135 1.425 ;
      RECT  8.285 1.425 9.13 1.43 ;
      RECT  8.285 1.43 9.125 1.435 ;
      RECT  8.285 1.435 9.12 1.44 ;
      RECT  8.285 1.44 9.115 1.445 ;
      RECT  8.285 1.445 9.11 1.45 ;
      RECT  8.285 1.45 9.105 1.455 ;
      RECT  8.285 1.455 9.1 1.46 ;
      RECT  8.285 1.46 9.095 1.465 ;
      RECT  8.285 1.465 9.09 1.47 ;
      RECT  8.285 1.47 9.085 1.475 ;
      RECT  8.285 1.475 9.08 1.48 ;
      RECT  8.285 1.48 9.075 1.485 ;
      RECT  8.285 1.485 9.07 1.49 ;
      RECT  8.285 1.49 9.065 1.495 ;
      RECT  8.285 1.495 9.06 1.5 ;
      RECT  8.285 1.5 9.055 1.505 ;
      RECT  8.285 1.505 9.05 1.51 ;
      RECT  8.285 1.51 9.045 1.515 ;
      RECT  8.285 1.515 9.04 1.52 ;
      RECT  8.285 1.52 9.035 1.525 ;
      RECT  8.285 1.525 9.03 1.53 ;
      RECT  8.285 1.53 9.025 1.535 ;
      RECT  8.285 1.535 9.02 1.54 ;
      RECT  8.285 1.54 9.015 1.545 ;
      RECT  8.285 1.545 9.01 1.55 ;
      RECT  8.285 1.55 9.005 1.555 ;
      RECT  8.285 1.555 9.0 1.56 ;
      RECT  8.285 1.56 8.995 1.565 ;
      RECT  8.285 1.565 8.99 1.57 ;
      RECT  8.285 1.57 8.985 1.575 ;
      RECT  8.285 1.575 8.98 1.58 ;
      RECT  8.285 1.58 8.515 1.81 ;
      RECT  5.43 1.75 5.77 1.81 ;
      RECT  5.43 1.81 8.515 2.04 ;
      RECT  6.605 2.04 6.835 3.245 ;
      RECT  5.43 3.245 7.24 3.475 ;
      RECT  17.19 0.37 17.53 0.6 ;
      RECT  17.19 0.6 17.42 1.005 ;
      RECT  14.445 0.37 16.355 0.6 ;
      RECT  16.125 0.6 16.355 1.005 ;
      RECT  14.445 0.6 14.675 1.35 ;
      RECT  16.125 1.005 17.42 1.235 ;
      RECT  9.965 1.29 12.45 1.35 ;
      RECT  9.965 1.35 14.675 1.52 ;
      RECT  12.18 1.52 14.675 1.58 ;
      RECT  9.965 1.52 10.195 3.315 ;
      RECT  4.015 0.83 6.54 1.06 ;
      RECT  6.2 1.06 6.54 1.12 ;
      RECT  4.015 1.06 4.245 1.29 ;
      RECT  9.47 0.83 13.26 1.06 ;
      RECT  12.92 1.06 13.26 1.12 ;
      RECT  9.47 1.06 9.7 1.75 ;
      RECT  9.14 1.75 9.7 1.98 ;
      RECT  7.49 0.89 8.78 1.12 ;
      RECT  7.49 1.12 7.72 1.35 ;
      RECT  4.66 1.29 6.005 1.295 ;
      RECT  4.66 1.295 6.01 1.3 ;
      RECT  4.66 1.3 6.015 1.305 ;
      RECT  4.66 1.305 6.02 1.31 ;
      RECT  4.66 1.31 6.025 1.315 ;
      RECT  4.66 1.315 6.03 1.32 ;
      RECT  4.66 1.32 6.035 1.325 ;
      RECT  4.66 1.325 6.04 1.33 ;
      RECT  4.66 1.33 6.045 1.335 ;
      RECT  4.66 1.335 6.05 1.34 ;
      RECT  4.66 1.34 6.055 1.345 ;
      RECT  4.66 1.345 6.06 1.35 ;
      RECT  4.66 1.35 7.72 1.52 ;
      RECT  5.9 1.52 7.72 1.525 ;
      RECT  4.66 1.52 5.0 1.56 ;
      RECT  5.905 1.525 7.72 1.53 ;
      RECT  5.91 1.53 7.72 1.535 ;
      RECT  5.915 1.535 7.72 1.54 ;
      RECT  5.92 1.54 7.72 1.545 ;
      RECT  5.925 1.545 7.72 1.55 ;
      RECT  5.93 1.55 7.72 1.555 ;
      RECT  5.935 1.555 7.72 1.56 ;
      RECT  5.94 1.56 7.72 1.565 ;
      RECT  5.945 1.565 7.72 1.57 ;
      RECT  5.95 1.57 7.72 1.575 ;
      RECT  5.955 1.575 7.72 1.58 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 1.81 ;
      RECT  12.82 1.81 15.235 2.04 ;
      RECT  12.82 2.04 13.05 2.335 ;
      RECT  15.005 2.04 15.235 2.38 ;
      RECT  12.71 2.335 13.05 2.565 ;
      RECT  15.005 2.38 16.41 2.61 ;
      RECT  15.005 2.61 15.235 3.805 ;
      RECT  13.62 3.805 15.5 4.035 ;
      RECT  10.68 1.75 11.72 1.98 ;
      RECT  11.085 1.98 11.315 3.545 ;
      RECT  8.285 2.35 8.515 3.245 ;
      RECT  8.285 3.245 9.7 3.475 ;
      RECT  9.47 3.475 9.7 3.545 ;
      RECT  9.47 3.545 11.72 3.775 ;
      RECT  8.77 2.66 9.15 2.685 ;
      RECT  8.77 2.685 9.635 2.915 ;
      RECT  9.405 2.35 9.635 2.685 ;
      RECT  8.77 2.915 9.15 2.94 ;
      RECT  5.97 2.355 6.35 2.94 ;
      RECT  3.96 4.215 5.0 4.445 ;
      RECT  6.2 4.215 8.78 4.445 ;
      RECT  0.18 4.365 1.85 4.595 ;
      RECT  1.51 4.595 1.85 4.675 ;
      RECT  1.51 4.675 8.475 4.905 ;
      RECT  8.245 4.905 8.475 5.0 ;
      RECT  1.51 4.905 1.85 5.23 ;
      RECT  4.87 4.905 5.21 5.23 ;
      RECT  8.245 5.0 10.81 5.23 ;
      RECT  10.68 4.48 13.26 4.71 ;
      LAYER METAL2 ;
      RECT  5.97 2.66 9.15 2.94 ;
      LAYER VIA12 ;
      RECT  6.03 2.67 6.29 2.93 ;
      RECT  8.83 2.67 9.09 2.93 ;
  END
END MDN_FDNRB_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNRB_2
#      Description : D-Flip Flop, neg-edge triggered, lo-async-clear
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNRB_2
  CLASS CORE ;
  FOREIGN MDN_FDNRB_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.86 1.565 17.74 1.795 ;
      RECT  16.685 1.795 16.915 3.245 ;
      RECT  15.86 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.1 1.565 19.98 1.795 ;
      RECT  18.925 1.795 19.155 3.245 ;
      RECT  18.1 3.245 19.98 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END QN
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.885 2.355 14.115 2.685 ;
      RECT  12.205 2.685 14.115 2.915 ;
      RECT  12.205 2.915 12.435 4.02 ;
      RECT  7.11 2.405 7.955 2.635 ;
      RECT  7.725 2.635 7.955 3.755 ;
      RECT  2.66 2.125 2.94 3.755 ;
      RECT  2.66 3.755 9.27 3.985 ;
      RECT  9.04 3.985 9.27 4.02 ;
      RECT  9.04 4.02 12.435 4.25 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  12.205 4.94 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 4.87 14.675 5.46 ;
      RECT  7.67 5.135 8.01 5.46 ;
      RECT  7.28 5.46 8.4 5.74 ;
      RECT  3.19 5.135 3.53 5.46 ;
      RECT  2.8 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  12.205 -0.14 14.115 0.14 ;
      RECT  12.205 0.14 12.435 0.6 ;
      RECT  13.885 0.14 14.115 0.89 ;
      RECT  13.62 0.89 14.115 1.12 ;
      RECT  6.72 -0.14 7.28 0.14 ;
      RECT  7.05 0.14 7.28 0.89 ;
      RECT  6.9 0.89 7.28 1.12 ;
      RECT  2.24 -0.14 2.915 0.14 ;
      RECT  2.685 0.14 2.915 1.005 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 1.74 1.235 ;
      RECT  3.24 0.37 6.33 0.6 ;
      RECT  3.24 0.6 3.47 1.565 ;
      RECT  1.565 1.565 3.47 1.795 ;
      RECT  1.565 1.795 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  9.01 0.37 11.93 0.6 ;
      RECT  9.01 0.6 9.24 1.225 ;
      RECT  9.005 1.225 9.24 1.23 ;
      RECT  9.0 1.23 9.24 1.235 ;
      RECT  8.995 1.235 9.24 1.24 ;
      RECT  8.99 1.24 9.24 1.245 ;
      RECT  8.985 1.245 9.24 1.25 ;
      RECT  8.98 1.25 9.24 1.255 ;
      RECT  8.975 1.255 9.24 1.26 ;
      RECT  8.97 1.26 9.24 1.265 ;
      RECT  8.965 1.265 9.24 1.27 ;
      RECT  8.96 1.27 9.24 1.275 ;
      RECT  8.955 1.275 9.24 1.28 ;
      RECT  8.95 1.28 9.24 1.285 ;
      RECT  8.945 1.285 9.24 1.29 ;
      RECT  8.94 1.29 9.24 1.295 ;
      RECT  8.935 1.295 9.24 1.3 ;
      RECT  8.93 1.3 9.24 1.305 ;
      RECT  8.925 1.305 9.24 1.31 ;
      RECT  8.92 1.31 9.24 1.315 ;
      RECT  8.915 1.315 9.24 1.32 ;
      RECT  8.91 1.32 9.235 1.325 ;
      RECT  8.905 1.325 9.23 1.33 ;
      RECT  8.9 1.33 9.225 1.335 ;
      RECT  8.895 1.335 9.22 1.34 ;
      RECT  8.89 1.34 9.215 1.345 ;
      RECT  8.885 1.345 9.21 1.35 ;
      RECT  8.285 1.35 9.205 1.355 ;
      RECT  8.285 1.355 9.2 1.36 ;
      RECT  8.285 1.36 9.195 1.365 ;
      RECT  8.285 1.365 9.19 1.37 ;
      RECT  8.285 1.37 9.185 1.375 ;
      RECT  8.285 1.375 9.18 1.38 ;
      RECT  8.285 1.38 9.175 1.385 ;
      RECT  8.285 1.385 9.17 1.39 ;
      RECT  8.285 1.39 9.165 1.395 ;
      RECT  8.285 1.395 9.16 1.4 ;
      RECT  8.285 1.4 9.155 1.405 ;
      RECT  8.285 1.405 9.15 1.41 ;
      RECT  8.285 1.41 9.145 1.415 ;
      RECT  8.285 1.415 9.14 1.42 ;
      RECT  8.285 1.42 9.135 1.425 ;
      RECT  8.285 1.425 9.13 1.43 ;
      RECT  8.285 1.43 9.125 1.435 ;
      RECT  8.285 1.435 9.12 1.44 ;
      RECT  8.285 1.44 9.115 1.445 ;
      RECT  8.285 1.445 9.11 1.45 ;
      RECT  8.285 1.45 9.105 1.455 ;
      RECT  8.285 1.455 9.1 1.46 ;
      RECT  8.285 1.46 9.095 1.465 ;
      RECT  8.285 1.465 9.09 1.47 ;
      RECT  8.285 1.47 9.085 1.475 ;
      RECT  8.285 1.475 9.08 1.48 ;
      RECT  8.285 1.48 9.075 1.485 ;
      RECT  8.285 1.485 9.07 1.49 ;
      RECT  8.285 1.49 9.065 1.495 ;
      RECT  8.285 1.495 9.06 1.5 ;
      RECT  8.285 1.5 9.055 1.505 ;
      RECT  8.285 1.505 9.05 1.51 ;
      RECT  8.285 1.51 9.045 1.515 ;
      RECT  8.285 1.515 9.04 1.52 ;
      RECT  8.285 1.52 9.035 1.525 ;
      RECT  8.285 1.525 9.03 1.53 ;
      RECT  8.285 1.53 9.025 1.535 ;
      RECT  8.285 1.535 9.02 1.54 ;
      RECT  8.285 1.54 9.015 1.545 ;
      RECT  8.285 1.545 9.01 1.55 ;
      RECT  8.285 1.55 9.005 1.555 ;
      RECT  8.285 1.555 9.0 1.56 ;
      RECT  8.285 1.56 8.995 1.565 ;
      RECT  8.285 1.565 8.99 1.57 ;
      RECT  8.285 1.57 8.985 1.575 ;
      RECT  8.285 1.575 8.98 1.58 ;
      RECT  8.285 1.58 8.515 1.81 ;
      RECT  5.43 1.75 5.77 1.81 ;
      RECT  5.43 1.81 8.515 2.04 ;
      RECT  6.605 2.04 6.835 3.245 ;
      RECT  5.43 3.245 7.24 3.475 ;
      RECT  19.43 0.37 19.77 0.6 ;
      RECT  19.43 0.6 19.66 1.005 ;
      RECT  18.31 0.37 18.65 0.6 ;
      RECT  18.42 0.6 18.65 1.005 ;
      RECT  14.445 0.37 16.355 0.6 ;
      RECT  16.125 0.6 16.355 1.005 ;
      RECT  14.445 0.6 14.675 1.565 ;
      RECT  16.125 1.005 19.66 1.235 ;
      RECT  10.015 1.29 12.435 1.52 ;
      RECT  12.205 1.52 12.435 1.565 ;
      RECT  10.015 1.52 10.245 3.315 ;
      RECT  12.205 1.565 14.675 1.795 ;
      RECT  3.96 0.83 6.54 1.06 ;
      RECT  6.2 1.06 6.54 1.12 ;
      RECT  3.96 1.06 4.3 1.205 ;
      RECT  9.47 0.83 13.26 1.06 ;
      RECT  12.92 1.06 13.26 1.12 ;
      RECT  9.47 1.06 9.7 1.75 ;
      RECT  9.14 1.75 9.7 1.98 ;
      RECT  7.725 0.89 8.78 1.12 ;
      RECT  7.725 1.12 7.955 1.35 ;
      RECT  4.66 1.29 6.01 1.295 ;
      RECT  4.66 1.295 6.015 1.3 ;
      RECT  4.66 1.3 6.02 1.305 ;
      RECT  4.66 1.305 6.025 1.31 ;
      RECT  4.66 1.31 6.03 1.315 ;
      RECT  4.66 1.315 6.035 1.32 ;
      RECT  4.66 1.32 6.04 1.325 ;
      RECT  4.66 1.325 6.045 1.33 ;
      RECT  4.66 1.33 6.05 1.335 ;
      RECT  4.66 1.335 6.055 1.34 ;
      RECT  4.66 1.34 6.06 1.345 ;
      RECT  4.66 1.345 6.065 1.35 ;
      RECT  4.66 1.35 7.955 1.52 ;
      RECT  5.905 1.52 7.955 1.525 ;
      RECT  5.91 1.525 7.955 1.53 ;
      RECT  5.915 1.53 7.955 1.535 ;
      RECT  5.92 1.535 7.955 1.54 ;
      RECT  5.925 1.54 7.955 1.545 ;
      RECT  5.93 1.545 7.955 1.55 ;
      RECT  5.935 1.55 7.955 1.555 ;
      RECT  5.94 1.555 7.955 1.56 ;
      RECT  5.945 1.56 7.955 1.565 ;
      RECT  5.95 1.565 7.955 1.57 ;
      RECT  5.955 1.57 7.955 1.575 ;
      RECT  5.96 1.575 7.955 1.58 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 4.365 ;
      RECT  13.62 4.365 17.42 4.595 ;
      RECT  13.62 4.595 13.85 5.0 ;
      RECT  16.18 4.595 16.41 5.0 ;
      RECT  17.19 4.595 17.42 5.0 ;
      RECT  12.71 5.0 13.85 5.23 ;
      RECT  16.07 5.0 16.41 5.23 ;
      RECT  17.19 5.0 17.53 5.23 ;
      RECT  10.525 1.75 11.72 1.98 ;
      RECT  10.525 1.98 10.755 3.245 ;
      RECT  10.525 3.245 11.72 3.475 ;
      RECT  10.525 3.475 10.755 3.55 ;
      RECT  8.285 2.35 8.515 3.245 ;
      RECT  8.285 3.245 9.785 3.475 ;
      RECT  9.555 3.475 9.785 3.55 ;
      RECT  9.555 3.55 10.755 3.775 ;
      RECT  9.555 3.775 10.735 3.78 ;
      RECT  5.97 2.355 6.35 2.94 ;
      RECT  9.33 2.365 9.71 2.94 ;
      RECT  3.96 4.215 4.595 4.365 ;
      RECT  3.96 4.365 5.0 4.445 ;
      RECT  4.365 4.445 5.0 4.595 ;
      RECT  6.2 4.215 8.78 4.445 ;
      RECT  10.68 4.48 13.26 4.71 ;
      RECT  7.165 4.675 8.515 4.905 ;
      RECT  7.165 4.905 7.395 5.0 ;
      RECT  8.285 4.905 8.515 5.0 ;
      RECT  0.18 4.365 1.85 4.595 ;
      RECT  1.51 4.595 1.85 4.675 ;
      RECT  1.51 4.675 4.035 4.905 ;
      RECT  3.805 4.905 4.035 5.0 ;
      RECT  1.51 4.905 1.85 5.23 ;
      RECT  3.805 5.0 7.395 5.23 ;
      RECT  8.285 5.0 10.81 5.23 ;
      LAYER METAL2 ;
      RECT  5.97 2.66 9.71 2.94 ;
      LAYER VIA12 ;
      RECT  6.03 2.67 6.29 2.93 ;
      RECT  9.39 2.67 9.65 2.93 ;
  END
END MDN_FDNRB_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNRBQ_F_1
#      Description : D-Flip Flop, neg-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNRBQ_F_1
  CLASS CORE ;
  FOREIGN MDN_FDNRBQ_F_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.98 0.37 1.85 0.6 ;
      RECT  0.98 0.6 1.26 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.245 1.565 17.74 1.795 ;
      RECT  17.245 1.795 17.475 3.245 ;
      RECT  17.245 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.885 4.41 15.18 4.64 ;
      RECT  13.885 4.64 14.115 4.925 ;
      RECT  14.95 4.64 15.18 5.0 ;
      RECT  7.165 4.41 10.755 4.64 ;
      RECT  7.165 4.64 7.395 4.925 ;
      RECT  10.525 4.64 10.755 4.925 ;
      RECT  8.23 4.64 8.57 5.23 ;
      RECT  0.42 4.36 2.355 4.41 ;
      RECT  0.42 4.41 3.935 4.59 ;
      RECT  2.125 4.59 3.935 4.64 ;
      RECT  0.42 4.59 0.7 5.0 ;
      RECT  3.705 4.64 3.935 4.925 ;
      RECT  3.705 4.925 7.395 5.155 ;
      RECT  10.525 4.925 14.115 5.155 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  14.95 5.0 15.29 5.23 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 10.64 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.56 -0.14 15.235 0.14 ;
      RECT  15.005 0.14 15.235 1.005 ;
      RECT  15.005 1.005 15.5 1.235 ;
      RECT  8.285 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.565 ;
      RECT  8.285 0.14 8.515 1.005 ;
      RECT  8.285 1.005 8.78 1.235 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 10.81 0.6 ;
      RECT  10.47 0.6 10.7 0.795 ;
      RECT  9.195 0.795 10.7 1.025 ;
      RECT  9.195 1.025 9.425 1.29 ;
      RECT  11.085 0.37 13.05 0.6 ;
      RECT  11.085 0.6 11.315 1.255 ;
      RECT  9.94 1.255 11.315 1.485 ;
      RECT  9.94 1.485 10.17 1.52 ;
      RECT  4.87 0.37 5.21 0.375 ;
      RECT  4.87 0.375 7.96 0.605 ;
      RECT  7.73 0.605 7.96 1.52 ;
      RECT  7.73 1.52 10.17 1.75 ;
      RECT  12.92 0.89 13.96 1.12 ;
      RECT  1.72 1.005 5.0 1.235 ;
      RECT  6.2 1.005 7.24 1.235 ;
      RECT  12.15 1.35 13.72 1.58 ;
      RECT  13.49 1.58 13.72 3.49 ;
      RECT  12.15 3.49 16.275 3.495 ;
      RECT  12.15 3.495 16.3 3.72 ;
      RECT  16.07 3.72 16.3 4.365 ;
      RECT  16.07 4.365 17.42 4.595 ;
      RECT  16.07 4.595 16.3 5.0 ;
      RECT  17.19 4.595 17.42 5.0 ;
      RECT  16.07 5.0 16.41 5.23 ;
      RECT  17.19 5.0 17.53 5.23 ;
      RECT  2.42 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 2.41 ;
      RECT  3.245 2.41 4.09 2.64 ;
      RECT  3.245 2.64 3.475 3.245 ;
      RECT  2.42 3.245 3.475 3.475 ;
      RECT  3.245 3.475 3.475 3.49 ;
      RECT  3.245 3.49 11.875 3.72 ;
      RECT  6.045 2.35 6.275 3.49 ;
      RECT  11.645 2.35 11.875 3.49 ;
      RECT  3.955 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 3.03 ;
      RECT  3.96 3.03 5.155 3.26 ;
      RECT  13.95 1.565 16.2 1.795 ;
      RECT  13.95 1.795 14.18 3.03 ;
      RECT  13.95 3.03 16.2 3.26 ;
      RECT  10.68 1.75 11.72 1.81 ;
      RECT  10.68 1.81 12.435 1.98 ;
      RECT  11.085 1.98 12.435 2.04 ;
      RECT  11.085 2.04 11.315 3.03 ;
      RECT  12.205 2.04 12.435 3.03 ;
      RECT  10.68 3.03 11.315 3.26 ;
      RECT  12.205 3.03 13.26 3.26 ;
      RECT  7.165 1.98 10.24 2.21 ;
      RECT  10.01 2.21 10.24 2.435 ;
      RECT  7.165 2.21 7.395 2.735 ;
      RECT  10.01 2.435 10.675 2.665 ;
      RECT  10.01 2.665 10.24 3.03 ;
      RECT  9.1 3.03 10.24 3.26 ;
      RECT  8.55 2.445 9.69 2.675 ;
      RECT  8.55 2.675 8.78 3.03 ;
      RECT  5.43 1.565 6.835 1.795 ;
      RECT  5.43 1.795 5.66 3.03 ;
      RECT  6.605 1.795 6.835 3.03 ;
      RECT  5.43 3.03 5.77 3.26 ;
      RECT  6.605 3.03 8.78 3.26 ;
      RECT  1.72 3.805 2.915 3.95 ;
      RECT  1.72 3.95 4.395 4.035 ;
      RECT  2.685 4.035 4.395 4.18 ;
      RECT  4.165 4.18 4.395 4.41 ;
      RECT  4.165 4.41 6.54 4.64 ;
      RECT  4.66 3.95 7.24 4.18 ;
      RECT  11.38 3.95 15.5 4.18 ;
  END
END MDN_FDNRBQ_F_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNRBQ_F_2
#      Description : D-Flip Flop, neg-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNRBQ_F_2
  CLASS CORE ;
  FOREIGN MDN_FDNRBQ_F_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.98 0.37 1.85 0.6 ;
      RECT  0.98 0.6 1.26 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.4 1.565 18.44 1.795 ;
      RECT  17.805 1.795 18.035 3.245 ;
      RECT  17.4 3.245 18.44 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.96 4.49 15.16 4.72 ;
      RECT  13.96 4.72 14.19 4.925 ;
      RECT  14.93 4.72 15.16 5.0 ;
      RECT  7.725 4.365 10.755 4.435 ;
      RECT  7.15 4.435 10.755 4.595 ;
      RECT  7.15 4.595 8.44 4.665 ;
      RECT  10.525 4.595 10.755 4.925 ;
      RECT  7.15 4.665 7.38 4.925 ;
      RECT  8.21 4.665 8.44 5.0 ;
      RECT  0.42 4.34 1.235 4.44 ;
      RECT  0.42 4.44 3.935 4.67 ;
      RECT  3.705 4.67 3.935 4.925 ;
      RECT  0.42 4.67 0.7 5.0 ;
      RECT  3.705 4.925 7.38 5.155 ;
      RECT  10.525 4.925 14.19 5.155 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  8.21 5.0 8.57 5.23 ;
      RECT  14.93 5.0 15.29 5.23 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.925 16.915 5.46 ;
      RECT  16.685 5.46 20.33 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  14.445 4.955 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  18.07 5.47 18.33 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.56 -0.14 15.235 0.14 ;
      RECT  15.005 0.14 15.235 1.005 ;
      RECT  15.005 1.005 15.5 1.235 ;
      RECT  8.285 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.565 ;
      RECT  8.285 0.14 8.515 1.005 ;
      RECT  8.285 1.005 8.78 1.235 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 10.81 0.6 ;
      RECT  10.47 0.6 10.7 0.795 ;
      RECT  9.195 0.795 10.7 1.025 ;
      RECT  9.195 1.025 9.425 1.29 ;
      RECT  11.085 0.37 13.05 0.6 ;
      RECT  11.085 0.6 11.315 1.255 ;
      RECT  9.94 1.255 11.315 1.485 ;
      RECT  9.94 1.485 10.17 1.525 ;
      RECT  4.87 0.37 5.21 0.445 ;
      RECT  4.87 0.445 7.96 0.675 ;
      RECT  7.73 0.675 7.96 1.525 ;
      RECT  7.73 1.525 10.17 1.755 ;
      RECT  12.92 0.96 13.96 1.19 ;
      RECT  1.72 1.005 5.0 1.235 ;
      RECT  6.2 1.005 7.24 1.235 ;
      RECT  12.15 1.42 13.775 1.65 ;
      RECT  13.545 1.65 13.775 3.56 ;
      RECT  12.15 3.56 16.3 3.79 ;
      RECT  16.07 3.79 16.3 4.365 ;
      RECT  16.07 4.365 17.42 4.595 ;
      RECT  16.07 4.595 16.3 5.0 ;
      RECT  17.19 4.595 17.42 5.0 ;
      RECT  16.07 5.0 16.41 5.23 ;
      RECT  17.19 5.0 18.65 5.23 ;
      RECT  2.42 1.565 3.47 1.795 ;
      RECT  3.24 1.795 3.47 2.405 ;
      RECT  3.24 2.405 4.09 2.635 ;
      RECT  3.24 2.635 3.47 3.515 ;
      RECT  2.42 3.515 11.875 3.745 ;
      RECT  6.045 2.35 6.275 3.515 ;
      RECT  11.645 2.35 11.875 3.515 ;
      RECT  3.955 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 3.055 ;
      RECT  3.96 3.055 5.155 3.285 ;
      RECT  14.075 1.565 16.2 1.795 ;
      RECT  14.075 1.795 14.305 3.1 ;
      RECT  14.075 3.1 16.2 3.33 ;
      RECT  10.68 1.715 11.72 1.88 ;
      RECT  10.68 1.88 12.955 1.945 ;
      RECT  11.09 1.945 12.955 2.11 ;
      RECT  11.09 2.11 11.32 3.055 ;
      RECT  12.725 2.11 12.955 3.1 ;
      RECT  10.68 3.055 11.32 3.285 ;
      RECT  12.725 3.1 13.26 3.33 ;
      RECT  7.165 1.985 10.195 2.215 ;
      RECT  9.965 2.215 10.195 2.4 ;
      RECT  7.165 2.215 7.395 2.69 ;
      RECT  9.965 2.4 10.81 2.63 ;
      RECT  9.965 2.63 10.195 3.055 ;
      RECT  9.14 3.055 10.195 3.285 ;
      RECT  8.55 2.445 9.69 2.675 ;
      RECT  8.55 2.675 8.78 3.055 ;
      RECT  5.43 1.75 6.835 1.98 ;
      RECT  5.43 1.98 5.66 3.055 ;
      RECT  6.605 1.98 6.835 3.055 ;
      RECT  5.43 3.055 5.77 3.285 ;
      RECT  6.605 3.055 8.78 3.285 ;
      RECT  1.72 3.975 4.4 4.205 ;
      RECT  4.17 4.205 4.4 4.465 ;
      RECT  4.17 4.465 6.54 4.695 ;
      RECT  4.66 3.975 7.27 4.205 ;
      RECT  11.38 4.025 15.5 4.255 ;
  END
END MDN_FDNRBQ_F_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNRBQ_F_4
#      Description : D-Flip Flop, neg-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNRBQ_F_4
  CLASS CORE ;
  FOREIGN MDN_FDNRBQ_F_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.98 0.37 1.85 0.6 ;
      RECT  0.98 0.6 1.26 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.4 1.565 20.68 1.795 ;
      RECT  20.045 1.795 20.275 3.245 ;
      RECT  17.4 3.245 20.685 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.97 4.415 15.18 4.645 ;
      RECT  13.97 4.645 14.2 4.925 ;
      RECT  14.95 4.645 15.18 5.0 ;
      RECT  7.15 4.425 10.715 4.655 ;
      RECT  7.15 4.655 7.38 4.925 ;
      RECT  10.485 4.655 10.715 4.925 ;
      RECT  8.23 4.655 8.46 5.0 ;
      RECT  0.42 4.34 1.235 4.425 ;
      RECT  0.42 4.425 3.935 4.655 ;
      RECT  3.705 4.655 3.935 4.925 ;
      RECT  0.42 4.655 0.7 5.0 ;
      RECT  3.705 4.925 7.38 5.155 ;
      RECT  10.485 4.925 14.2 5.155 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  8.23 5.0 8.57 5.23 ;
      RECT  14.95 5.0 15.29 5.23 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 22.57 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  9.965 4.93 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  20.31 5.47 20.57 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.925 -0.14 19.6 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.56 -0.14 15.235 0.14 ;
      RECT  15.005 0.14 15.235 1.005 ;
      RECT  15.005 1.005 15.5 1.235 ;
      RECT  8.285 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.6 ;
      RECT  8.285 0.14 8.515 1.005 ;
      RECT  8.285 1.005 8.78 1.235 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 10.81 0.6 ;
      RECT  10.47 0.6 10.7 0.83 ;
      RECT  9.195 0.83 10.7 1.06 ;
      RECT  9.195 1.06 9.425 1.29 ;
      RECT  11.085 0.37 13.05 0.6 ;
      RECT  11.085 0.6 11.315 1.29 ;
      RECT  9.965 1.29 11.315 1.52 ;
      RECT  9.965 1.52 10.195 1.525 ;
      RECT  4.87 0.37 5.21 0.445 ;
      RECT  4.87 0.445 7.955 0.675 ;
      RECT  7.725 0.675 7.955 1.525 ;
      RECT  7.725 1.525 10.195 1.755 ;
      RECT  1.72 1.005 5.0 1.235 ;
      RECT  6.2 1.005 7.24 1.235 ;
      RECT  12.92 1.005 13.96 1.235 ;
      RECT  3.955 1.565 5.095 1.795 ;
      RECT  4.865 1.795 5.095 2.35 ;
      RECT  4.865 2.35 5.1 2.69 ;
      RECT  4.865 2.69 5.095 3.03 ;
      RECT  3.96 3.03 5.095 3.26 ;
      RECT  13.95 1.565 16.2 1.795 ;
      RECT  13.95 1.795 14.18 3.035 ;
      RECT  13.95 3.035 16.2 3.265 ;
      RECT  10.68 1.75 11.72 1.93 ;
      RECT  10.68 1.93 12.955 1.98 ;
      RECT  11.085 1.98 12.955 2.16 ;
      RECT  11.085 2.16 11.315 3.03 ;
      RECT  12.725 2.16 12.955 3.035 ;
      RECT  10.68 3.03 11.315 3.26 ;
      RECT  12.725 3.035 13.26 3.265 ;
      RECT  7.165 1.985 10.24 2.215 ;
      RECT  10.01 2.215 10.24 2.4 ;
      RECT  7.165 2.215 7.395 2.69 ;
      RECT  10.01 2.4 10.81 2.63 ;
      RECT  10.01 2.63 10.24 3.03 ;
      RECT  9.1 3.03 10.24 3.26 ;
      RECT  16.07 2.405 19.675 2.635 ;
      RECT  16.685 2.635 16.915 3.495 ;
      RECT  12.15 1.465 13.72 1.695 ;
      RECT  13.49 1.695 13.72 3.495 ;
      RECT  12.15 3.495 16.915 3.725 ;
      RECT  11.645 2.41 11.985 2.64 ;
      RECT  11.645 2.64 11.875 3.49 ;
      RECT  2.42 1.565 3.45 1.795 ;
      RECT  3.22 1.795 3.45 2.405 ;
      RECT  3.22 2.405 4.09 2.635 ;
      RECT  3.22 2.635 3.45 3.49 ;
      RECT  2.42 3.49 11.875 3.72 ;
      RECT  6.045 2.35 6.275 3.49 ;
      RECT  8.55 2.445 9.69 2.675 ;
      RECT  8.55 2.675 8.78 3.03 ;
      RECT  5.43 1.75 6.835 1.98 ;
      RECT  5.43 1.98 5.66 3.03 ;
      RECT  6.605 1.98 6.835 3.03 ;
      RECT  5.43 3.03 5.77 3.26 ;
      RECT  6.605 3.03 8.78 3.26 ;
      RECT  1.72 3.95 4.395 4.18 ;
      RECT  4.165 4.18 4.395 4.465 ;
      RECT  4.165 4.465 6.54 4.695 ;
      RECT  4.66 3.95 7.24 4.18 ;
      RECT  11.38 3.955 15.5 4.185 ;
      RECT  19.43 5.0 20.89 5.23 ;
  END
END MDN_FDNRBQ_F_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNRBQ_1
#      Description : D-Flip Flop, neg-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNRBQ_1
  CLASS CORE ;
  FOREIGN MDN_FDNRBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 3.245 ;
      RECT  15.005 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 9.66 2.355 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  9.965 4.925 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 4.925 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  8.4 -0.14 9.52 0.14 ;
      RECT  8.845 0.14 9.075 0.89 ;
      RECT  8.44 0.89 9.48 1.12 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.6 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  12.7 0.37 13.04 0.375 ;
      RECT  9.94 0.375 13.04 0.6 ;
      RECT  9.94 0.6 12.955 0.605 ;
      RECT  9.94 0.605 10.17 1.39 ;
      RECT  4.87 0.37 5.21 0.83 ;
      RECT  1.775 0.83 5.69 1.005 ;
      RECT  1.775 1.005 7.93 1.06 ;
      RECT  5.46 1.06 7.93 1.235 ;
      RECT  1.775 1.06 2.005 1.565 ;
      RECT  7.7 1.235 7.93 1.39 ;
      RECT  7.7 1.39 10.17 1.62 ;
      RECT  1.565 1.565 2.005 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 2.06 4.035 ;
      RECT  14.95 0.37 15.29 0.6 ;
      RECT  14.95 0.6 15.18 1.005 ;
      RECT  10.68 1.005 15.18 1.235 ;
      RECT  14.445 1.235 14.675 2.35 ;
      RECT  13.885 2.35 14.675 2.58 ;
      RECT  13.885 2.58 14.115 4.005 ;
      RECT  9.105 4.005 14.115 4.225 ;
      RECT  9.105 4.225 14.1 4.235 ;
      RECT  2.42 1.29 5.0 1.52 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  12.15 1.565 12.49 1.795 ;
      RECT  12.205 1.795 12.435 2.405 ;
      RECT  10.47 2.405 12.435 2.635 ;
      RECT  12.205 2.635 12.435 3.085 ;
      RECT  12.15 3.085 12.49 3.315 ;
      RECT  12.92 1.565 13.96 1.795 ;
      RECT  11.435 1.63 11.665 1.905 ;
      RECT  9.965 1.905 11.665 2.135 ;
      RECT  9.965 2.135 10.195 3.545 ;
      RECT  3.245 1.75 4.3 1.98 ;
      RECT  3.245 1.98 3.475 3.545 ;
      RECT  3.245 3.545 13.26 3.775 ;
      RECT  7.165 2.35 7.395 3.545 ;
      RECT  5.485 1.625 5.715 2.405 ;
      RECT  3.75 2.405 5.715 2.635 ;
      RECT  5.485 2.635 5.715 3.315 ;
      RECT  2.42 4.005 6.54 4.235 ;
      RECT  6.77 4.005 8.78 4.235 ;
      RECT  6.77 4.235 7.0 4.465 ;
      RECT  4.66 4.465 7.0 4.695 ;
      RECT  7.23 4.465 10.755 4.695 ;
      RECT  7.23 4.695 7.46 5.0 ;
      RECT  10.525 4.695 10.755 5.0 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.465 ;
      RECT  0.18 4.465 3.995 4.695 ;
      RECT  3.765 4.695 3.995 5.0 ;
      RECT  1.51 4.695 1.85 5.23 ;
      RECT  3.765 5.0 7.46 5.23 ;
      RECT  10.525 5.0 11.93 5.23 ;
      RECT  11.38 4.475 13.96 4.705 ;
  END
END MDN_FDNRBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNRBQ_2
#      Description : D-Flip Flop, neg-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNRBQ_2
  CLASS CORE ;
  FOREIGN MDN_FDNRBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.16 1.565 16.2 1.795 ;
      RECT  15.565 1.795 15.795 3.245 ;
      RECT  15.16 3.245 16.2 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 9.66 2.355 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  9.965 4.925 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 4.925 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.245 4.93 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.925 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  8.4 -0.14 9.52 0.14 ;
      RECT  8.845 0.14 9.075 1.005 ;
      RECT  8.44 1.005 9.48 1.235 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.6 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  9.97 0.37 13.05 0.6 ;
      RECT  9.97 0.6 10.2 1.465 ;
      RECT  4.87 0.37 5.21 0.83 ;
      RECT  1.775 0.83 5.69 1.005 ;
      RECT  1.775 1.005 7.955 1.06 ;
      RECT  5.46 1.06 7.955 1.235 ;
      RECT  1.775 1.06 2.005 1.565 ;
      RECT  7.725 1.235 7.955 1.465 ;
      RECT  7.725 1.465 10.205 1.695 ;
      RECT  1.565 1.565 2.005 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 2.06 4.035 ;
      RECT  14.95 0.37 16.41 0.6 ;
      RECT  10.68 1.005 14.675 1.235 ;
      RECT  14.445 1.235 14.675 2.405 ;
      RECT  13.83 2.405 15.23 2.635 ;
      RECT  13.885 2.635 14.115 4.005 ;
      RECT  9.105 4.005 14.115 4.235 ;
      RECT  2.42 1.29 5.0 1.52 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  12.92 1.565 13.96 1.795 ;
      RECT  11.435 1.51 11.665 1.94 ;
      RECT  9.965 1.94 11.665 2.17 ;
      RECT  9.965 2.17 10.195 3.545 ;
      RECT  3.245 1.75 4.3 1.98 ;
      RECT  3.245 1.98 3.475 3.545 ;
      RECT  3.245 3.545 13.26 3.775 ;
      RECT  7.165 2.35 7.395 3.545 ;
      RECT  5.485 1.51 5.715 2.405 ;
      RECT  3.75 2.405 5.715 2.635 ;
      RECT  5.485 2.635 5.715 3.315 ;
      RECT  12.205 1.51 12.435 2.405 ;
      RECT  10.47 2.405 12.435 2.635 ;
      RECT  12.205 2.635 12.435 3.315 ;
      RECT  2.475 3.75 2.705 4.005 ;
      RECT  2.475 4.005 6.54 4.235 ;
      RECT  6.805 4.005 8.78 4.235 ;
      RECT  6.805 4.235 7.035 4.48 ;
      RECT  4.66 4.48 7.035 4.71 ;
      RECT  7.265 4.465 10.755 4.695 ;
      RECT  7.265 4.695 7.495 5.0 ;
      RECT  10.525 4.695 10.755 5.0 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.465 ;
      RECT  0.235 4.31 0.465 4.465 ;
      RECT  0.235 4.465 4.035 4.695 ;
      RECT  3.805 4.695 4.035 5.0 ;
      RECT  1.51 4.695 1.85 5.23 ;
      RECT  3.8 5.0 7.495 5.23 ;
      RECT  10.525 5.0 11.93 5.23 ;
      RECT  11.38 4.48 13.96 4.71 ;
  END
END MDN_FDNRBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNRBQ_4
#      Description : D-Flip Flop, neg-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNRBQ_4
  CLASS CORE ;
  FOREIGN MDN_FDNRBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.16 1.565 18.445 1.795 ;
      RECT  17.805 1.795 18.035 3.245 ;
      RECT  15.16 3.245 18.44 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 9.66 2.355 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  7.725 4.925 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 4.925 10.195 5.46 ;
      RECT  3.245 4.94 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.94 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  8.4 -0.14 9.52 0.14 ;
      RECT  8.845 0.14 9.075 1.005 ;
      RECT  8.44 1.005 9.48 1.235 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.6 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  9.965 0.37 13.05 0.6 ;
      RECT  9.965 0.6 10.195 1.485 ;
      RECT  4.87 0.37 5.21 0.83 ;
      RECT  1.775 0.83 5.715 1.005 ;
      RECT  1.775 1.005 7.955 1.06 ;
      RECT  5.485 1.06 7.955 1.235 ;
      RECT  1.775 1.06 2.005 1.565 ;
      RECT  7.725 1.235 7.955 1.485 ;
      RECT  7.725 1.485 10.195 1.715 ;
      RECT  1.565 1.565 2.005 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 2.06 4.035 ;
      RECT  17.18 0.37 18.65 0.6 ;
      RECT  10.68 1.005 14.675 1.235 ;
      RECT  14.445 1.235 14.675 2.405 ;
      RECT  13.83 2.405 17.325 2.635 ;
      RECT  13.885 2.635 14.115 4.005 ;
      RECT  9.105 4.005 14.115 4.235 ;
      RECT  2.475 1.29 5.0 1.52 ;
      RECT  2.475 1.52 2.705 1.85 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  12.92 1.565 13.96 1.795 ;
      RECT  11.435 1.51 11.665 1.945 ;
      RECT  9.965 1.945 11.665 2.175 ;
      RECT  9.965 2.175 10.195 3.545 ;
      RECT  3.245 1.75 4.3 1.98 ;
      RECT  3.245 1.98 3.475 3.545 ;
      RECT  3.245 3.545 13.26 3.775 ;
      RECT  7.165 2.35 7.395 3.545 ;
      RECT  5.485 1.51 5.715 2.405 ;
      RECT  3.75 2.405 5.715 2.635 ;
      RECT  5.485 2.635 5.715 3.315 ;
      RECT  12.205 1.51 12.435 2.405 ;
      RECT  10.47 2.405 12.435 2.635 ;
      RECT  12.205 2.635 12.435 3.315 ;
      RECT  2.42 4.005 6.54 4.235 ;
      RECT  6.77 4.005 8.78 4.235 ;
      RECT  6.77 4.235 7.0 4.48 ;
      RECT  4.66 4.48 7.0 4.71 ;
      RECT  7.26 4.465 10.755 4.695 ;
      RECT  7.26 4.695 7.49 5.0 ;
      RECT  10.525 4.695 10.755 5.0 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 1.74 4.48 ;
      RECT  0.18 4.48 4.035 4.595 ;
      RECT  1.51 4.595 4.035 4.71 ;
      RECT  1.51 4.71 1.74 5.0 ;
      RECT  3.805 4.71 4.035 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  3.805 5.0 7.49 5.23 ;
      RECT  10.525 5.0 11.93 5.23 ;
      RECT  11.38 4.48 13.96 4.71 ;
  END
END MDN_FDNRBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNRBSBQ_1
#      Description : D-Flip Flop neg-edge triggered, lo-async-clear/set, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNRBSBQ_1
  CLASS CORE ;
  FOREIGN MDN_FDNRBSBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  2.42 3.245 2.915 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 1.565 11.9 2.125 ;
      RECT  8.285 2.125 11.9 2.355 ;
      RECT  8.285 2.355 8.515 2.69 ;
      RECT  11.62 2.355 11.9 2.69 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.47 0.37 16.915 0.6 ;
      RECT  16.685 0.6 16.915 1.565 ;
      RECT  16.685 1.565 17.5 1.795 ;
      RECT  17.22 1.795 17.5 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  12.205 5.08 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.965 5.08 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 5.08 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.245 5.0 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  17.245 -0.14 18.09 0.14 ;
      RECT  17.245 0.14 17.475 1.005 ;
      RECT  17.245 1.005 17.74 1.235 ;
      RECT  9.52 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 1.005 ;
      RECT  8.44 1.005 11.72 1.235 ;
      RECT  2.8 -0.14 3.92 0.14 ;
      RECT  3.19 0.14 3.53 0.51 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  4.925 0.37 6.33 0.6 ;
      RECT  4.925 0.6 5.155 0.74 ;
      RECT  3.245 0.74 5.155 0.97 ;
      RECT  3.245 0.97 3.475 1.005 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 3.475 1.235 ;
      RECT  7.725 0.37 9.69 0.6 ;
      RECT  7.725 0.6 7.955 1.005 ;
      RECT  5.485 1.005 7.955 1.235 ;
      RECT  5.485 1.235 5.715 3.39 ;
      RECT  13.62 1.005 16.2 1.235 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  12.205 1.565 13.26 1.795 ;
      RECT  12.205 1.795 12.435 3.24 ;
      RECT  11.38 3.24 13.26 3.47 ;
      RECT  13.885 1.565 14.73 1.795 ;
      RECT  13.885 1.795 14.115 2.415 ;
      RECT  12.71 2.415 14.115 2.645 ;
      RECT  13.885 2.645 14.115 3.24 ;
      RECT  13.885 3.24 14.73 3.47 ;
      RECT  15.16 1.565 16.355 1.795 ;
      RECT  16.125 1.795 16.355 3.7 ;
      RECT  7.725 1.565 9.48 1.795 ;
      RECT  7.725 1.795 7.955 2.025 ;
      RECT  7.165 2.025 7.955 2.255 ;
      RECT  7.165 2.255 7.395 3.16 ;
      RECT  7.165 3.16 9.635 3.39 ;
      RECT  9.405 3.39 9.635 3.7 ;
      RECT  9.405 3.7 16.355 3.93 ;
      RECT  6.045 2.35 6.275 2.66 ;
      RECT  6.045 2.66 6.91 2.94 ;
      RECT  15.005 2.345 15.235 2.66 ;
      RECT  14.37 2.66 15.235 2.94 ;
      RECT  4.925 2.35 5.155 3.16 ;
      RECT  3.805 3.16 5.155 3.245 ;
      RECT  3.245 3.245 5.155 3.39 ;
      RECT  3.245 3.39 4.035 3.475 ;
      RECT  3.245 3.475 3.475 3.805 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 3.475 4.035 ;
      RECT  4.66 3.62 8.78 3.85 ;
      RECT  3.96 4.08 6.54 4.31 ;
      RECT  6.77 4.16 14.675 4.39 ;
      RECT  6.77 4.39 7.0 4.54 ;
      RECT  14.445 4.39 14.675 5.0 ;
      RECT  2.74 4.54 7.0 4.77 ;
      RECT  2.74 4.77 2.97 5.0 ;
      RECT  2.63 5.0 2.97 5.23 ;
      RECT  14.445 5.0 16.41 5.23 ;
      RECT  0.18 4.365 1.74 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  15.16 4.365 17.74 4.595 ;
      RECT  7.23 4.62 14.06 4.85 ;
      RECT  7.23 4.85 7.46 5.0 ;
      RECT  13.83 4.85 14.06 5.0 ;
      RECT  4.87 5.0 7.46 5.23 ;
      RECT  13.83 5.0 14.17 5.23 ;
      LAYER METAL2 ;
      RECT  6.53 2.66 14.75 2.94 ;
      LAYER VIA12 ;
      RECT  6.59 2.67 6.85 2.93 ;
      RECT  14.43 2.67 14.69 2.93 ;
  END
END MDN_FDNRBSBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNRBSBQ_2
#      Description : D-Flip Flop neg-edge triggered, lo-async-clear/set, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNRBSBQ_2
  CLASS CORE ;
  FOREIGN MDN_FDNRBSBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.1 1.565 19.98 1.795 ;
      RECT  18.925 1.795 19.155 3.245 ;
      RECT  18.1 3.245 19.98 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.285 2.125 11.9 2.355 ;
      RECT  8.285 2.355 8.515 2.69 ;
      RECT  11.62 2.355 11.9 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.22 4.365 17.5 5.0 ;
      RECT  17.19 5.0 17.53 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  12.15 5.085 12.49 5.46 ;
      RECT  11.76 5.46 12.88 5.74 ;
      RECT  7.67 5.085 8.01 5.46 ;
      RECT  7.28 5.46 10.64 5.74 ;
      RECT  9.91 5.085 10.25 5.46 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  17.36 -0.14 18.48 0.14 ;
      RECT  17.805 0.14 18.035 1.005 ;
      RECT  17.4 1.005 18.035 1.235 ;
      RECT  8.4 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 1.005 ;
      RECT  8.44 1.005 11.72 1.235 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.52 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  18.07 -0.13 18.33 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.445 ;
      RECT  3.705 0.445 6.33 0.675 ;
      RECT  3.705 0.675 3.935 0.75 ;
      RECT  2.63 0.37 2.97 0.75 ;
      RECT  1.565 0.75 3.935 0.98 ;
      RECT  1.565 0.98 1.795 1.565 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  7.725 0.37 9.69 0.6 ;
      RECT  7.725 0.6 7.955 1.005 ;
      RECT  5.485 1.005 7.955 1.235 ;
      RECT  5.485 1.235 5.715 3.53 ;
      RECT  10.47 0.37 17.53 0.6 ;
      RECT  19.43 0.37 19.77 0.6 ;
      RECT  19.43 0.6 19.66 1.005 ;
      RECT  18.31 0.37 18.65 0.6 ;
      RECT  18.42 0.6 18.65 1.005 ;
      RECT  18.42 1.005 19.66 1.235 ;
      RECT  13.03 0.83 16.915 1.06 ;
      RECT  13.03 1.06 13.26 1.565 ;
      RECT  16.685 1.06 16.915 2.405 ;
      RECT  12.205 1.565 13.26 1.795 ;
      RECT  12.205 1.795 12.435 3.245 ;
      RECT  16.07 2.405 18.65 2.635 ;
      RECT  11.38 3.245 13.26 3.475 ;
      RECT  13.62 1.29 16.2 1.52 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  2.42 1.665 2.915 1.895 ;
      RECT  2.685 1.895 2.915 3.245 ;
      RECT  2.42 3.245 5.155 3.475 ;
      RECT  4.925 2.35 5.155 3.245 ;
      RECT  13.885 1.75 14.73 1.98 ;
      RECT  13.885 1.98 14.115 2.415 ;
      RECT  12.71 2.415 14.115 2.645 ;
      RECT  13.885 2.645 14.115 3.245 ;
      RECT  13.885 3.245 14.73 3.475 ;
      RECT  15.005 1.75 15.5 1.98 ;
      RECT  15.005 1.98 15.235 3.705 ;
      RECT  7.725 1.565 9.48 1.795 ;
      RECT  7.725 1.795 7.955 2.405 ;
      RECT  7.11 2.405 7.955 2.635 ;
      RECT  7.725 2.635 7.955 3.145 ;
      RECT  7.725 3.145 10.195 3.375 ;
      RECT  9.965 3.375 10.195 3.705 ;
      RECT  9.965 3.705 15.235 3.935 ;
      RECT  6.045 2.35 6.275 3.245 ;
      RECT  6.045 3.245 7.45 3.475 ;
      RECT  7.22 3.475 7.45 3.605 ;
      RECT  7.22 3.605 9.62 3.835 ;
      RECT  9.39 3.835 9.62 4.165 ;
      RECT  9.39 4.165 14.675 4.395 ;
      RECT  14.445 4.395 14.675 5.0 ;
      RECT  14.445 5.0 15.29 5.23 ;
      RECT  15.565 3.245 17.74 3.475 ;
      RECT  15.565 3.475 15.795 4.365 ;
      RECT  15.16 4.365 15.795 4.595 ;
      RECT  4.66 3.805 6.99 4.035 ;
      RECT  6.76 4.035 6.99 4.065 ;
      RECT  6.76 4.065 8.78 4.295 ;
      RECT  3.96 4.365 6.54 4.595 ;
      RECT  7.165 4.625 14.06 4.855 ;
      RECT  7.165 4.855 7.395 5.0 ;
      RECT  13.83 4.855 14.06 5.0 ;
      RECT  4.87 5.0 7.395 5.23 ;
      RECT  13.83 5.0 14.17 5.23 ;
  END
END MDN_FDNRBSBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNRBSBQ_4
#      Description : D-Flip Flop neg-edge triggered, lo-async-clear/set, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNRBSBQ_4
  CLASS CORE ;
  FOREIGN MDN_FDNRBSBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.805 1.565 22.22 1.795 ;
      RECT  20.045 1.795 20.275 3.245 ;
      RECT  18.09 3.245 22.22 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.845 2.115 11.875 2.125 ;
      RECT  8.845 2.125 11.9 2.345 ;
      RECT  8.845 2.345 9.075 2.38 ;
      RECT  11.62 2.345 11.9 2.915 ;
      RECT  8.77 2.38 9.075 2.405 ;
      RECT  8.23 2.405 9.075 2.635 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.22 4.365 17.5 5.0 ;
      RECT  17.19 5.0 17.53 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.905 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.905 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.905 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 12.88 5.74 ;
      RECT  12.15 5.135 12.49 5.46 ;
      RECT  7.67 5.135 8.01 5.46 ;
      RECT  7.28 5.46 8.4 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.695 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 1.005 ;
      RECT  17.4 1.005 19.155 1.235 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 1.005 ;
      RECT  8.44 1.005 11.72 1.235 ;
      RECT  2.8 -0.14 3.92 0.14 ;
      RECT  3.19 0.14 3.53 0.465 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  9.35 0.37 9.69 0.375 ;
      RECT  7.725 0.375 9.69 0.6 ;
      RECT  7.725 0.6 9.645 0.605 ;
      RECT  7.725 0.605 7.955 1.445 ;
      RECT  5.485 1.445 7.955 1.675 ;
      RECT  5.485 1.675 5.715 3.53 ;
      RECT  5.485 0.37 6.33 0.6 ;
      RECT  5.485 0.6 5.715 0.695 ;
      RECT  2.62 0.37 2.96 0.695 ;
      RECT  1.775 0.695 5.715 0.925 ;
      RECT  1.775 0.925 2.005 3.455 ;
      RECT  10.47 0.37 17.53 0.6 ;
      RECT  13.03 0.83 16.915 1.06 ;
      RECT  13.03 1.06 13.26 1.565 ;
      RECT  16.685 1.06 16.915 2.405 ;
      RECT  12.205 1.565 13.26 1.795 ;
      RECT  12.205 1.795 12.435 3.245 ;
      RECT  16.07 2.405 19.675 2.635 ;
      RECT  11.38 3.245 13.26 3.475 ;
      RECT  6.2 0.89 7.24 1.12 ;
      RECT  3.915 1.155 5.0 1.385 ;
      RECT  13.62 1.29 16.2 1.52 ;
      RECT  2.475 1.615 5.155 1.845 ;
      RECT  4.925 1.845 5.155 2.69 ;
      RECT  2.475 1.845 2.705 3.475 ;
      RECT  14.39 1.75 14.73 1.98 ;
      RECT  14.42 1.98 14.7 2.685 ;
      RECT  12.765 2.35 12.995 2.685 ;
      RECT  12.765 2.685 14.7 2.915 ;
      RECT  14.42 2.915 14.7 3.46 ;
      RECT  15.005 1.75 15.5 1.98 ;
      RECT  15.005 1.98 15.235 3.755 ;
      RECT  8.285 1.565 9.48 1.795 ;
      RECT  8.285 1.795 8.515 1.94 ;
      RECT  7.165 1.94 8.515 2.17 ;
      RECT  7.165 2.17 7.395 3.03 ;
      RECT  7.165 3.03 10.195 3.26 ;
      RECT  9.965 3.26 10.195 3.755 ;
      RECT  9.965 3.755 15.235 3.985 ;
      RECT  20.55 2.405 22.01 2.635 ;
      RECT  15.565 3.245 17.74 3.475 ;
      RECT  15.565 3.475 15.795 4.365 ;
      RECT  15.11 4.365 15.795 4.595 ;
      RECT  6.045 2.35 6.275 3.56 ;
      RECT  6.045 3.56 9.635 3.79 ;
      RECT  9.405 3.79 9.635 4.215 ;
      RECT  9.405 4.215 14.675 4.445 ;
      RECT  14.445 4.445 14.675 5.0 ;
      RECT  14.445 5.0 15.29 5.23 ;
      RECT  4.64 4.02 8.78 4.25 ;
      RECT  3.96 4.48 6.54 4.71 ;
      RECT  7.165 4.675 14.06 4.905 ;
      RECT  7.165 4.905 7.395 5.0 ;
      RECT  13.83 4.905 14.06 5.0 ;
      RECT  4.87 5.0 7.395 5.23 ;
      RECT  13.83 5.0 14.17 5.23 ;
      RECT  19.43 5.0 20.89 5.23 ;
  END
END MDN_FDNRBSBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNSBQ_1
#      Description : D-Flip Flop neg-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNSBQ_1
  CLASS CORE ;
  FOREIGN MDN_FDNSBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 3.245 ;
      RECT  15.005 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.57 1.565 13.02 1.795 ;
      RECT  11.57 1.795 11.875 1.945 ;
      RECT  12.74 1.795 13.02 2.915 ;
      RECT  8.285 1.945 11.875 2.175 ;
      RECT  8.285 2.175 8.515 2.69 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.87 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  7.725 5.075 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 5.08 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 1.005 ;
      RECT  12.92 1.005 14.675 1.235 ;
      RECT  8.285 -0.14 8.96 0.14 ;
      RECT  8.285 0.14 8.515 1.005 ;
      RECT  8.285 1.005 8.78 1.235 ;
      RECT  5.04 -0.14 6.16 0.14 ;
      RECT  5.43 0.14 5.77 0.465 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  13.83 0.37 14.17 0.445 ;
      RECT  9.91 0.445 14.17 0.675 ;
      RECT  3.245 0.44 3.475 0.695 ;
      RECT  3.245 0.695 7.45 0.925 ;
      RECT  7.11 0.37 7.45 0.695 ;
      RECT  9.14 1.005 11.72 1.235 ;
      RECT  2.42 1.155 6.54 1.385 ;
      RECT  6.9 1.485 11.02 1.715 ;
      RECT  6.9 1.715 7.13 2.405 ;
      RECT  6.17 2.405 7.13 2.635 ;
      RECT  6.9 2.635 7.13 3.155 ;
      RECT  6.9 3.155 9.48 3.385 ;
      RECT  13.62 1.565 14.115 1.795 ;
      RECT  13.885 1.795 14.115 3.245 ;
      RECT  11.535 2.445 11.875 2.675 ;
      RECT  11.645 2.675 11.875 3.245 ;
      RECT  11.645 3.245 14.115 3.475 ;
      RECT  13.885 3.475 14.115 4.365 ;
      RECT  13.885 4.365 15.18 4.595 ;
      RECT  14.95 4.595 15.18 5.0 ;
      RECT  14.95 5.0 15.29 5.23 ;
      RECT  3.96 1.615 5.0 1.845 ;
      RECT  9.35 2.405 10.195 2.635 ;
      RECT  9.965 2.635 10.195 3.615 ;
      RECT  3.805 2.355 4.035 3.215 ;
      RECT  3.805 3.215 6.275 3.32 ;
      RECT  3.8 3.32 6.275 3.325 ;
      RECT  3.795 3.325 6.275 3.33 ;
      RECT  3.79 3.33 6.275 3.335 ;
      RECT  3.785 3.335 6.275 3.34 ;
      RECT  3.78 3.34 6.275 3.345 ;
      RECT  3.775 3.345 6.275 3.35 ;
      RECT  3.77 3.35 6.275 3.355 ;
      RECT  3.765 3.355 6.275 3.36 ;
      RECT  3.76 3.36 6.275 3.365 ;
      RECT  3.755 3.365 6.275 3.37 ;
      RECT  3.75 3.37 6.275 3.375 ;
      RECT  3.745 3.375 6.275 3.38 ;
      RECT  3.74 3.38 6.275 3.385 ;
      RECT  3.735 3.385 6.275 3.39 ;
      RECT  3.73 3.39 6.275 3.395 ;
      RECT  3.725 3.395 6.275 3.4 ;
      RECT  3.72 3.4 6.275 3.405 ;
      RECT  3.715 3.405 6.275 3.41 ;
      RECT  3.71 3.41 6.275 3.415 ;
      RECT  3.705 3.415 6.275 3.42 ;
      RECT  3.7 3.42 6.275 3.425 ;
      RECT  3.695 3.425 6.275 3.43 ;
      RECT  3.69 3.43 6.275 3.435 ;
      RECT  3.685 3.435 6.275 3.44 ;
      RECT  3.68 3.44 6.275 3.445 ;
      RECT  3.675 3.445 4.0 3.45 ;
      RECT  6.045 3.445 6.275 3.615 ;
      RECT  3.67 3.45 3.995 3.455 ;
      RECT  3.665 3.455 3.99 3.46 ;
      RECT  3.66 3.46 3.985 3.465 ;
      RECT  3.655 3.465 3.98 3.47 ;
      RECT  3.65 3.47 3.975 3.475 ;
      RECT  3.645 3.475 3.97 3.48 ;
      RECT  3.64 3.48 3.965 3.485 ;
      RECT  3.635 3.485 3.96 3.49 ;
      RECT  3.63 3.49 3.955 3.495 ;
      RECT  3.625 3.495 3.95 3.5 ;
      RECT  3.62 3.5 3.945 3.505 ;
      RECT  3.615 3.505 3.94 3.51 ;
      RECT  3.61 3.51 3.935 3.515 ;
      RECT  3.605 3.515 3.93 3.52 ;
      RECT  3.6 3.52 3.925 3.525 ;
      RECT  3.595 3.525 3.92 3.53 ;
      RECT  3.59 3.53 3.915 3.535 ;
      RECT  3.585 3.535 3.91 3.54 ;
      RECT  3.58 3.54 3.905 3.545 ;
      RECT  3.575 3.545 3.9 3.55 ;
      RECT  3.57 3.55 3.895 3.555 ;
      RECT  3.565 3.555 3.89 3.56 ;
      RECT  3.56 3.56 3.885 3.565 ;
      RECT  3.555 3.565 3.88 3.57 ;
      RECT  3.55 3.57 3.875 3.575 ;
      RECT  3.545 3.575 3.87 3.58 ;
      RECT  3.54 3.58 3.865 3.585 ;
      RECT  3.535 3.585 3.86 3.59 ;
      RECT  3.53 3.59 3.855 3.595 ;
      RECT  3.525 3.595 3.85 3.6 ;
      RECT  3.52 3.6 3.845 3.605 ;
      RECT  3.515 3.605 3.84 3.61 ;
      RECT  3.51 3.61 3.835 3.615 ;
      RECT  3.505 3.615 3.83 3.62 ;
      RECT  6.045 3.615 10.195 3.845 ;
      RECT  3.5 3.62 3.825 3.625 ;
      RECT  3.495 3.625 3.82 3.63 ;
      RECT  3.49 3.63 3.815 3.635 ;
      RECT  3.485 3.635 3.81 3.64 ;
      RECT  3.48 3.64 3.805 3.645 ;
      RECT  3.475 3.645 3.8 3.65 ;
      RECT  3.47 3.65 3.795 3.655 ;
      RECT  3.465 3.655 3.79 3.66 ;
      RECT  3.46 3.66 3.785 3.665 ;
      RECT  3.455 3.665 3.78 3.67 ;
      RECT  3.45 3.67 3.775 3.675 ;
      RECT  3.445 3.675 3.77 3.68 ;
      RECT  3.44 3.68 3.765 3.685 ;
      RECT  3.435 3.685 3.76 3.69 ;
      RECT  3.43 3.69 3.755 3.695 ;
      RECT  3.425 3.695 3.75 3.7 ;
      RECT  3.42 3.7 3.745 3.705 ;
      RECT  3.415 3.705 3.74 3.71 ;
      RECT  3.41 3.71 3.735 3.715 ;
      RECT  3.405 3.715 3.73 3.72 ;
      RECT  3.4 3.72 3.725 3.725 ;
      RECT  3.395 3.725 3.72 3.73 ;
      RECT  3.39 3.73 3.715 3.735 ;
      RECT  3.385 3.735 3.71 3.74 ;
      RECT  3.38 3.74 3.705 3.745 ;
      RECT  3.375 3.745 3.7 3.75 ;
      RECT  3.37 3.75 3.695 3.755 ;
      RECT  3.365 3.755 3.69 3.76 ;
      RECT  3.36 3.76 3.685 3.765 ;
      RECT  3.355 3.765 3.68 3.77 ;
      RECT  3.35 3.77 3.675 3.775 ;
      RECT  3.345 3.775 3.67 3.78 ;
      RECT  3.34 3.78 3.665 3.785 ;
      RECT  3.335 3.785 3.66 3.79 ;
      RECT  3.33 3.79 3.655 3.795 ;
      RECT  3.325 3.795 3.65 3.8 ;
      RECT  3.32 3.8 3.645 3.805 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 3.64 3.81 ;
      RECT  1.565 3.81 3.635 3.815 ;
      RECT  1.565 3.815 3.63 3.82 ;
      RECT  1.565 3.82 3.625 3.825 ;
      RECT  1.565 3.825 3.62 3.83 ;
      RECT  1.565 3.83 3.615 3.835 ;
      RECT  1.565 3.835 3.61 3.84 ;
      RECT  1.565 3.84 3.605 3.845 ;
      RECT  1.565 3.845 3.6 3.85 ;
      RECT  1.565 3.85 3.595 3.855 ;
      RECT  1.565 3.855 3.59 3.86 ;
      RECT  1.565 3.86 3.585 3.865 ;
      RECT  1.565 3.865 3.58 3.87 ;
      RECT  1.565 3.87 3.575 3.875 ;
      RECT  1.565 3.875 3.57 3.88 ;
      RECT  1.565 3.88 3.565 3.885 ;
      RECT  1.565 3.885 3.56 3.89 ;
      RECT  1.565 3.89 3.555 3.895 ;
      RECT  1.565 3.895 3.55 3.9 ;
      RECT  1.565 3.9 3.545 3.905 ;
      RECT  1.565 3.905 3.54 3.91 ;
      RECT  1.565 3.91 3.535 3.915 ;
      RECT  1.565 3.915 3.53 3.92 ;
      RECT  1.565 3.92 3.525 3.925 ;
      RECT  1.565 3.925 3.52 3.93 ;
      RECT  1.565 3.93 3.515 3.935 ;
      RECT  1.565 3.935 3.51 3.94 ;
      RECT  1.565 3.94 3.505 3.945 ;
      RECT  1.565 3.945 3.5 3.95 ;
      RECT  1.565 3.95 3.495 3.955 ;
      RECT  1.565 3.955 3.49 3.96 ;
      RECT  1.565 3.96 3.485 3.965 ;
      RECT  1.565 3.965 3.48 3.97 ;
      RECT  1.565 3.97 3.475 3.975 ;
      RECT  1.565 3.975 3.47 3.98 ;
      RECT  1.565 3.98 3.465 3.985 ;
      RECT  1.565 3.985 3.46 3.99 ;
      RECT  1.565 3.99 3.455 3.995 ;
      RECT  1.565 3.995 3.45 4.0 ;
      RECT  1.565 4.0 3.445 4.005 ;
      RECT  1.565 4.005 3.44 4.01 ;
      RECT  1.565 4.01 3.435 4.015 ;
      RECT  1.565 4.015 3.43 4.02 ;
      RECT  1.565 4.02 3.425 4.025 ;
      RECT  1.565 4.025 3.42 4.03 ;
      RECT  1.565 4.03 3.415 4.035 ;
      RECT  3.245 1.615 3.475 3.315 ;
      RECT  4.105 3.675 5.715 3.905 ;
      RECT  5.485 3.905 5.715 4.075 ;
      RECT  4.105 3.905 4.335 4.08 ;
      RECT  5.485 4.075 6.54 4.305 ;
      RECT  3.96 4.08 4.335 4.31 ;
      RECT  10.68 3.805 13.26 4.035 ;
      RECT  4.565 4.135 5.0 4.365 ;
      RECT  4.565 4.365 4.795 4.54 ;
      RECT  2.475 4.31 2.705 4.54 ;
      RECT  2.475 4.54 4.795 4.77 ;
      RECT  9.91 4.365 13.0 4.595 ;
      RECT  12.77 4.595 13.0 5.0 ;
      RECT  12.77 5.0 14.17 5.23 ;
      RECT  5.025 4.615 8.515 4.845 ;
      RECT  5.025 4.845 5.255 5.0 ;
      RECT  8.285 4.845 8.515 5.0 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 1.74 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 5.255 5.23 ;
      RECT  8.285 5.0 10.81 5.23 ;
  END
END MDN_FDNSBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNSBQ_2
#      Description : D-Flip Flop neg-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNSBQ_2
  CLASS CORE ;
  FOREIGN MDN_FDNSBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.16 1.565 16.2 1.795 ;
      RECT  15.565 1.795 15.795 3.245 ;
      RECT  15.16 3.245 16.2 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 1.93 13.02 2.16 ;
      RECT  8.26 2.16 8.54 2.915 ;
      RECT  12.74 2.16 13.02 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  7.725 5.08 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 5.08 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.445 0.14 14.675 1.005 ;
      RECT  12.92 1.005 14.73 1.235 ;
      RECT  8.285 -0.14 8.96 0.14 ;
      RECT  8.285 0.14 8.515 1.005 ;
      RECT  8.285 1.005 8.78 1.235 ;
      RECT  5.04 -0.14 6.16 0.14 ;
      RECT  5.43 0.14 5.77 0.465 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 1.74 1.235 ;
      RECT  9.91 0.37 14.17 0.6 ;
      RECT  14.95 0.37 16.41 0.6 ;
      RECT  3.19 0.445 5.155 0.675 ;
      RECT  4.925 0.675 5.155 0.695 ;
      RECT  4.925 0.695 7.45 0.925 ;
      RECT  7.11 0.37 7.45 0.695 ;
      RECT  2.42 1.005 4.595 1.155 ;
      RECT  2.42 1.155 6.54 1.235 ;
      RECT  4.365 1.235 6.54 1.385 ;
      RECT  9.14 1.005 11.72 1.235 ;
      RECT  6.9 1.47 11.02 1.7 ;
      RECT  6.9 1.7 7.13 2.405 ;
      RECT  5.99 2.405 7.13 2.635 ;
      RECT  6.9 2.635 7.13 3.24 ;
      RECT  6.9 3.24 8.515 3.245 ;
      RECT  6.9 3.245 9.48 3.47 ;
      RECT  8.285 3.47 9.48 3.475 ;
      RECT  13.62 1.565 14.675 1.795 ;
      RECT  14.445 1.795 14.675 2.405 ;
      RECT  14.445 2.405 15.29 2.635 ;
      RECT  14.445 2.635 14.675 3.245 ;
      RECT  11.645 2.39 11.875 3.245 ;
      RECT  11.645 3.245 14.675 3.475 ;
      RECT  3.96 1.615 5.0 1.845 ;
      RECT  9.35 2.445 10.195 2.675 ;
      RECT  9.965 2.675 10.195 3.705 ;
      RECT  3.805 2.35 4.035 3.18 ;
      RECT  3.805 3.18 6.235 3.32 ;
      RECT  3.8 3.32 6.235 3.325 ;
      RECT  3.795 3.325 6.235 3.33 ;
      RECT  3.79 3.33 6.235 3.335 ;
      RECT  3.785 3.335 6.235 3.34 ;
      RECT  3.78 3.34 6.235 3.345 ;
      RECT  3.775 3.345 6.235 3.35 ;
      RECT  3.77 3.35 6.235 3.355 ;
      RECT  3.765 3.355 6.235 3.36 ;
      RECT  3.76 3.36 6.235 3.365 ;
      RECT  3.755 3.365 6.235 3.37 ;
      RECT  3.75 3.37 6.235 3.375 ;
      RECT  3.745 3.375 6.235 3.38 ;
      RECT  3.74 3.38 6.235 3.385 ;
      RECT  3.735 3.385 6.235 3.39 ;
      RECT  3.73 3.39 6.235 3.395 ;
      RECT  3.725 3.395 6.235 3.4 ;
      RECT  3.72 3.4 6.235 3.405 ;
      RECT  3.715 3.405 6.235 3.41 ;
      RECT  3.71 3.41 4.035 3.415 ;
      RECT  6.005 3.41 6.235 3.7 ;
      RECT  3.705 3.415 4.03 3.42 ;
      RECT  3.7 3.42 4.025 3.425 ;
      RECT  3.695 3.425 4.02 3.43 ;
      RECT  3.69 3.43 4.015 3.435 ;
      RECT  3.685 3.435 4.01 3.44 ;
      RECT  3.68 3.44 4.005 3.445 ;
      RECT  3.675 3.445 4.0 3.45 ;
      RECT  3.67 3.45 3.995 3.455 ;
      RECT  3.665 3.455 3.99 3.46 ;
      RECT  3.66 3.46 3.985 3.465 ;
      RECT  3.655 3.465 3.98 3.47 ;
      RECT  3.65 3.47 3.975 3.475 ;
      RECT  3.645 3.475 3.97 3.48 ;
      RECT  3.64 3.48 3.965 3.485 ;
      RECT  3.635 3.485 3.96 3.49 ;
      RECT  3.63 3.49 3.955 3.495 ;
      RECT  3.625 3.495 3.95 3.5 ;
      RECT  3.62 3.5 3.945 3.505 ;
      RECT  3.615 3.505 3.94 3.51 ;
      RECT  3.61 3.51 3.935 3.515 ;
      RECT  3.605 3.515 3.93 3.52 ;
      RECT  3.6 3.52 3.925 3.525 ;
      RECT  3.595 3.525 3.92 3.53 ;
      RECT  3.59 3.53 3.915 3.535 ;
      RECT  3.585 3.535 3.91 3.54 ;
      RECT  3.58 3.54 3.905 3.545 ;
      RECT  3.575 3.545 3.9 3.55 ;
      RECT  3.57 3.55 3.895 3.555 ;
      RECT  3.565 3.555 3.89 3.56 ;
      RECT  3.56 3.56 3.885 3.565 ;
      RECT  3.555 3.565 3.88 3.57 ;
      RECT  3.55 3.57 3.875 3.575 ;
      RECT  3.545 3.575 3.87 3.58 ;
      RECT  3.54 3.58 3.865 3.585 ;
      RECT  3.535 3.585 3.86 3.59 ;
      RECT  3.53 3.59 3.855 3.595 ;
      RECT  3.525 3.595 3.85 3.6 ;
      RECT  3.52 3.6 3.845 3.605 ;
      RECT  3.515 3.605 3.84 3.61 ;
      RECT  3.51 3.61 3.835 3.615 ;
      RECT  3.505 3.615 3.83 3.62 ;
      RECT  3.5 3.62 3.825 3.625 ;
      RECT  3.495 3.625 3.82 3.63 ;
      RECT  3.49 3.63 3.815 3.635 ;
      RECT  3.485 3.635 3.81 3.64 ;
      RECT  3.48 3.64 3.805 3.645 ;
      RECT  3.475 3.645 3.8 3.65 ;
      RECT  3.47 3.65 3.795 3.655 ;
      RECT  3.465 3.655 3.79 3.66 ;
      RECT  3.46 3.66 3.785 3.665 ;
      RECT  3.455 3.665 3.78 3.67 ;
      RECT  3.45 3.67 3.775 3.675 ;
      RECT  3.445 3.675 3.77 3.68 ;
      RECT  3.44 3.68 3.765 3.685 ;
      RECT  3.435 3.685 3.76 3.69 ;
      RECT  3.43 3.69 3.755 3.695 ;
      RECT  3.425 3.695 3.75 3.7 ;
      RECT  3.42 3.7 3.745 3.705 ;
      RECT  6.005 3.7 7.955 3.705 ;
      RECT  3.415 3.705 3.74 3.71 ;
      RECT  6.005 3.705 10.195 3.93 ;
      RECT  3.41 3.71 3.735 3.715 ;
      RECT  3.405 3.715 3.73 3.72 ;
      RECT  3.4 3.72 3.725 3.725 ;
      RECT  3.395 3.725 3.72 3.73 ;
      RECT  3.39 3.73 3.715 3.735 ;
      RECT  3.385 3.735 3.71 3.74 ;
      RECT  3.38 3.74 3.705 3.745 ;
      RECT  3.375 3.745 3.7 3.75 ;
      RECT  3.37 3.75 3.695 3.755 ;
      RECT  3.365 3.755 3.69 3.76 ;
      RECT  3.36 3.76 3.685 3.765 ;
      RECT  3.355 3.765 3.68 3.77 ;
      RECT  3.35 3.77 3.675 3.775 ;
      RECT  3.345 3.775 3.67 3.78 ;
      RECT  3.34 3.78 3.665 3.785 ;
      RECT  3.335 3.785 3.66 3.79 ;
      RECT  3.33 3.79 3.655 3.795 ;
      RECT  3.325 3.795 3.65 3.8 ;
      RECT  3.32 3.8 3.645 3.805 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.805 ;
      RECT  1.72 3.805 3.64 3.81 ;
      RECT  1.72 3.81 3.635 3.815 ;
      RECT  1.72 3.815 3.63 3.82 ;
      RECT  1.72 3.82 3.625 3.825 ;
      RECT  1.72 3.825 3.62 3.83 ;
      RECT  1.72 3.83 3.615 3.835 ;
      RECT  1.72 3.835 3.61 3.84 ;
      RECT  1.72 3.84 3.605 3.845 ;
      RECT  1.72 3.845 3.6 3.85 ;
      RECT  1.72 3.85 3.595 3.855 ;
      RECT  1.72 3.855 3.59 3.86 ;
      RECT  1.72 3.86 3.585 3.865 ;
      RECT  1.72 3.865 3.58 3.87 ;
      RECT  1.72 3.87 3.575 3.875 ;
      RECT  1.72 3.875 3.57 3.88 ;
      RECT  1.72 3.88 3.565 3.885 ;
      RECT  1.72 3.885 3.56 3.89 ;
      RECT  1.72 3.89 3.555 3.895 ;
      RECT  1.72 3.895 3.55 3.9 ;
      RECT  1.72 3.9 3.545 3.905 ;
      RECT  1.72 3.905 3.54 3.91 ;
      RECT  1.72 3.91 3.535 3.915 ;
      RECT  1.72 3.915 3.53 3.92 ;
      RECT  1.72 3.92 3.525 3.925 ;
      RECT  1.72 3.925 3.52 3.93 ;
      RECT  1.72 3.93 3.515 3.935 ;
      RECT  7.725 3.93 10.195 3.935 ;
      RECT  1.72 3.935 3.51 3.94 ;
      RECT  1.72 3.94 3.505 3.945 ;
      RECT  1.72 3.945 3.5 3.95 ;
      RECT  1.72 3.95 3.495 3.955 ;
      RECT  1.72 3.955 3.49 3.96 ;
      RECT  1.72 3.96 3.485 3.965 ;
      RECT  1.72 3.965 3.48 3.97 ;
      RECT  1.72 3.97 3.475 3.975 ;
      RECT  1.72 3.975 3.47 3.98 ;
      RECT  1.72 3.98 3.465 3.985 ;
      RECT  1.72 3.985 3.46 3.99 ;
      RECT  1.72 3.99 3.455 3.995 ;
      RECT  1.72 3.995 3.45 4.0 ;
      RECT  1.72 4.0 3.445 4.005 ;
      RECT  1.72 4.005 3.44 4.01 ;
      RECT  1.72 4.01 3.435 4.015 ;
      RECT  1.72 4.015 3.43 4.02 ;
      RECT  1.72 4.02 3.425 4.025 ;
      RECT  1.72 4.025 3.42 4.03 ;
      RECT  1.72 4.03 3.415 4.035 ;
      RECT  3.245 1.615 3.475 3.315 ;
      RECT  4.105 3.695 5.715 3.925 ;
      RECT  4.105 3.925 4.335 4.08 ;
      RECT  5.485 3.925 5.715 4.16 ;
      RECT  3.96 4.08 4.335 4.31 ;
      RECT  5.485 4.16 6.54 4.39 ;
      RECT  10.68 3.805 13.26 4.035 ;
      RECT  4.565 4.155 5.0 4.385 ;
      RECT  4.565 4.385 4.795 4.54 ;
      RECT  2.475 4.31 2.705 4.54 ;
      RECT  2.475 4.54 4.795 4.77 ;
      RECT  9.91 4.365 12.995 4.595 ;
      RECT  12.765 4.595 12.995 5.0 ;
      RECT  12.765 5.0 14.17 5.23 ;
      RECT  5.025 4.62 8.515 4.85 ;
      RECT  5.025 4.85 5.255 5.0 ;
      RECT  8.285 4.85 8.515 5.0 ;
      RECT  0.18 4.365 1.74 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 5.255 5.23 ;
      RECT  8.285 5.0 10.81 5.23 ;
  END
END MDN_FDNSBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FDNSBQ_4
#      Description : D-Flip Flop neg-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDNSBQ_4
  CLASS CORE ;
  FOREIGN MDN_FDNSBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.16 1.565 18.44 1.795 ;
      RECT  17.805 1.795 18.035 3.245 ;
      RECT  15.16 3.245 18.44 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.255 1.895 13.02 2.125 ;
      RECT  8.26 2.125 8.54 2.915 ;
      RECT  12.74 2.125 13.02 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  7.67 5.13 8.01 5.46 ;
      RECT  7.28 5.46 8.4 5.74 ;
      RECT  5.43 5.135 5.77 5.46 ;
      RECT  5.04 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 20.33 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  12.88 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 1.005 ;
      RECT  12.92 1.005 14.675 1.235 ;
      RECT  8.285 -0.14 8.96 0.14 ;
      RECT  8.285 0.14 8.515 0.97 ;
      RECT  8.285 0.97 8.78 1.2 ;
      RECT  5.04 -0.14 6.16 0.14 ;
      RECT  5.43 0.14 5.77 0.465 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  18.07 -0.13 18.33 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 1.74 1.235 ;
      RECT  7.11 0.37 7.45 0.6 ;
      RECT  7.11 0.6 7.34 0.695 ;
      RECT  3.19 0.445 5.155 0.675 ;
      RECT  4.925 0.675 5.155 0.695 ;
      RECT  4.925 0.695 7.34 0.925 ;
      RECT  9.91 0.37 14.17 0.6 ;
      RECT  17.19 0.37 18.65 0.6 ;
      RECT  2.42 1.005 4.595 1.16 ;
      RECT  2.42 1.16 6.54 1.235 ;
      RECT  4.365 1.235 6.54 1.39 ;
      RECT  9.14 0.965 11.72 1.195 ;
      RECT  6.77 1.435 11.02 1.665 ;
      RECT  6.77 1.665 7.0 2.405 ;
      RECT  6.135 2.405 7.0 2.635 ;
      RECT  6.77 2.635 7.0 3.245 ;
      RECT  6.77 3.245 9.48 3.475 ;
      RECT  8.44 3.24 8.78 3.245 ;
      RECT  13.62 1.565 14.675 1.795 ;
      RECT  14.445 1.795 14.675 2.405 ;
      RECT  14.445 2.405 17.435 2.635 ;
      RECT  14.445 2.635 14.675 3.245 ;
      RECT  11.645 2.355 11.875 3.245 ;
      RECT  11.645 3.245 14.675 3.475 ;
      RECT  3.96 1.62 5.0 1.85 ;
      RECT  9.35 2.435 9.945 2.665 ;
      RECT  9.715 2.665 9.945 3.74 ;
      RECT  3.805 2.34 4.035 3.245 ;
      RECT  3.805 3.245 6.275 3.32 ;
      RECT  6.045 3.24 6.275 3.245 ;
      RECT  3.8 3.32 6.275 3.325 ;
      RECT  3.795 3.325 6.275 3.33 ;
      RECT  3.79 3.33 6.275 3.335 ;
      RECT  3.785 3.335 6.275 3.34 ;
      RECT  3.78 3.34 6.275 3.345 ;
      RECT  3.775 3.345 6.275 3.35 ;
      RECT  3.77 3.35 6.275 3.355 ;
      RECT  3.765 3.355 6.275 3.36 ;
      RECT  3.76 3.36 6.275 3.365 ;
      RECT  3.755 3.365 6.275 3.37 ;
      RECT  3.75 3.37 6.275 3.375 ;
      RECT  3.745 3.375 6.275 3.38 ;
      RECT  3.74 3.38 6.275 3.385 ;
      RECT  3.735 3.385 6.275 3.39 ;
      RECT  3.73 3.39 6.275 3.395 ;
      RECT  3.725 3.395 6.275 3.4 ;
      RECT  3.72 3.4 6.275 3.405 ;
      RECT  3.715 3.405 6.275 3.41 ;
      RECT  3.71 3.41 6.275 3.415 ;
      RECT  3.705 3.415 6.275 3.42 ;
      RECT  3.7 3.42 6.275 3.425 ;
      RECT  3.695 3.425 6.275 3.43 ;
      RECT  3.69 3.43 6.275 3.435 ;
      RECT  3.685 3.435 6.275 3.44 ;
      RECT  3.68 3.44 6.275 3.445 ;
      RECT  3.675 3.445 6.275 3.45 ;
      RECT  3.67 3.45 6.275 3.455 ;
      RECT  3.665 3.455 6.275 3.46 ;
      RECT  3.66 3.46 6.275 3.465 ;
      RECT  3.655 3.465 6.275 3.47 ;
      RECT  3.65 3.47 6.275 3.475 ;
      RECT  3.645 3.475 3.97 3.48 ;
      RECT  6.045 3.475 6.275 3.74 ;
      RECT  3.64 3.48 3.965 3.485 ;
      RECT  3.635 3.485 3.96 3.49 ;
      RECT  3.63 3.49 3.955 3.495 ;
      RECT  3.625 3.495 3.95 3.5 ;
      RECT  3.62 3.5 3.945 3.505 ;
      RECT  3.615 3.505 3.94 3.51 ;
      RECT  3.61 3.51 3.935 3.515 ;
      RECT  3.605 3.515 3.93 3.52 ;
      RECT  3.6 3.52 3.925 3.525 ;
      RECT  3.595 3.525 3.92 3.53 ;
      RECT  3.59 3.53 3.915 3.535 ;
      RECT  3.585 3.535 3.91 3.54 ;
      RECT  3.58 3.54 3.905 3.545 ;
      RECT  3.575 3.545 3.9 3.55 ;
      RECT  3.57 3.55 3.895 3.555 ;
      RECT  3.565 3.555 3.89 3.56 ;
      RECT  3.56 3.56 3.885 3.565 ;
      RECT  3.555 3.565 3.88 3.57 ;
      RECT  3.55 3.57 3.875 3.575 ;
      RECT  3.545 3.575 3.87 3.58 ;
      RECT  3.54 3.58 3.865 3.585 ;
      RECT  3.535 3.585 3.86 3.59 ;
      RECT  3.53 3.59 3.855 3.595 ;
      RECT  3.525 3.595 3.85 3.6 ;
      RECT  3.52 3.6 3.845 3.605 ;
      RECT  3.515 3.605 3.84 3.61 ;
      RECT  3.51 3.61 3.835 3.615 ;
      RECT  3.505 3.615 3.83 3.62 ;
      RECT  3.5 3.62 3.825 3.625 ;
      RECT  3.495 3.625 3.82 3.63 ;
      RECT  3.49 3.63 3.815 3.635 ;
      RECT  3.485 3.635 3.81 3.64 ;
      RECT  3.48 3.64 3.805 3.645 ;
      RECT  3.475 3.645 3.8 3.65 ;
      RECT  3.47 3.65 3.795 3.655 ;
      RECT  3.465 3.655 3.79 3.66 ;
      RECT  3.46 3.66 3.785 3.665 ;
      RECT  3.455 3.665 3.78 3.67 ;
      RECT  3.45 3.67 3.775 3.675 ;
      RECT  3.445 3.675 3.77 3.68 ;
      RECT  3.44 3.68 3.765 3.685 ;
      RECT  3.435 3.685 3.76 3.69 ;
      RECT  3.43 3.69 3.755 3.695 ;
      RECT  3.425 3.695 3.75 3.7 ;
      RECT  3.42 3.7 3.745 3.705 ;
      RECT  3.415 3.705 3.74 3.71 ;
      RECT  3.41 3.71 3.735 3.715 ;
      RECT  3.405 3.715 3.73 3.72 ;
      RECT  3.4 3.72 3.725 3.725 ;
      RECT  3.395 3.725 3.72 3.73 ;
      RECT  3.39 3.73 3.715 3.735 ;
      RECT  3.385 3.735 3.71 3.74 ;
      RECT  3.38 3.74 3.705 3.745 ;
      RECT  6.045 3.74 9.945 3.97 ;
      RECT  3.375 3.745 3.7 3.75 ;
      RECT  3.37 3.75 3.695 3.755 ;
      RECT  3.365 3.755 3.69 3.76 ;
      RECT  3.36 3.76 3.685 3.765 ;
      RECT  3.355 3.765 3.68 3.77 ;
      RECT  3.35 3.77 3.675 3.775 ;
      RECT  3.345 3.775 3.67 3.78 ;
      RECT  3.34 3.78 3.665 3.785 ;
      RECT  3.335 3.785 3.66 3.79 ;
      RECT  3.33 3.79 3.655 3.795 ;
      RECT  3.325 3.795 3.65 3.8 ;
      RECT  3.32 3.8 3.645 3.805 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.805 ;
      RECT  1.72 3.805 3.64 3.81 ;
      RECT  1.72 3.81 3.635 3.815 ;
      RECT  1.72 3.815 3.63 3.82 ;
      RECT  1.72 3.82 3.625 3.825 ;
      RECT  1.72 3.825 3.62 3.83 ;
      RECT  1.72 3.83 3.615 3.835 ;
      RECT  1.72 3.835 3.61 3.84 ;
      RECT  1.72 3.84 3.605 3.845 ;
      RECT  1.72 3.845 3.6 3.85 ;
      RECT  1.72 3.85 3.595 3.855 ;
      RECT  1.72 3.855 3.59 3.86 ;
      RECT  1.72 3.86 3.585 3.865 ;
      RECT  1.72 3.865 3.58 3.87 ;
      RECT  1.72 3.87 3.575 3.875 ;
      RECT  1.72 3.875 3.57 3.88 ;
      RECT  1.72 3.88 3.565 3.885 ;
      RECT  1.72 3.885 3.56 3.89 ;
      RECT  1.72 3.89 3.555 3.895 ;
      RECT  1.72 3.895 3.55 3.9 ;
      RECT  1.72 3.9 3.545 3.905 ;
      RECT  1.72 3.905 3.54 3.91 ;
      RECT  1.72 3.91 3.535 3.915 ;
      RECT  1.72 3.915 3.53 3.92 ;
      RECT  1.72 3.92 3.525 3.925 ;
      RECT  1.72 3.925 3.52 3.93 ;
      RECT  1.72 3.93 3.515 3.935 ;
      RECT  1.72 3.935 3.51 3.94 ;
      RECT  1.72 3.94 3.505 3.945 ;
      RECT  1.72 3.945 3.5 3.95 ;
      RECT  1.72 3.95 3.495 3.955 ;
      RECT  1.72 3.955 3.49 3.96 ;
      RECT  1.72 3.96 3.485 3.965 ;
      RECT  1.72 3.965 3.48 3.97 ;
      RECT  1.72 3.97 3.475 3.975 ;
      RECT  1.72 3.975 3.47 3.98 ;
      RECT  1.72 3.98 3.465 3.985 ;
      RECT  1.72 3.985 3.46 3.99 ;
      RECT  1.72 3.99 3.455 3.995 ;
      RECT  1.72 3.995 3.45 4.0 ;
      RECT  1.72 4.0 3.445 4.005 ;
      RECT  1.72 4.005 3.44 4.01 ;
      RECT  1.72 4.01 3.435 4.015 ;
      RECT  1.72 4.015 3.43 4.02 ;
      RECT  1.72 4.02 3.425 4.025 ;
      RECT  1.72 4.025 3.42 4.03 ;
      RECT  1.72 4.03 3.415 4.035 ;
      RECT  3.245 1.62 3.475 3.315 ;
      RECT  10.68 3.805 13.26 4.035 ;
      RECT  3.96 3.85 5.715 4.08 ;
      RECT  5.485 4.08 5.715 4.205 ;
      RECT  5.485 4.205 6.54 4.435 ;
      RECT  2.42 4.31 5.0 4.54 ;
      RECT  9.91 4.365 12.995 4.595 ;
      RECT  12.765 4.595 12.995 5.0 ;
      RECT  12.765 5.0 14.17 5.23 ;
      RECT  5.24 4.665 8.515 4.67 ;
      RECT  5.235 4.67 8.515 4.675 ;
      RECT  5.23 4.675 8.515 4.68 ;
      RECT  5.225 4.68 8.515 4.685 ;
      RECT  5.22 4.685 8.515 4.69 ;
      RECT  5.215 4.69 8.515 4.695 ;
      RECT  5.21 4.695 8.515 4.7 ;
      RECT  5.205 4.7 8.515 4.705 ;
      RECT  5.2 4.705 8.515 4.71 ;
      RECT  5.195 4.71 8.515 4.715 ;
      RECT  5.19 4.715 8.515 4.72 ;
      RECT  5.185 4.72 8.515 4.725 ;
      RECT  5.18 4.725 8.515 4.73 ;
      RECT  5.175 4.73 8.515 4.735 ;
      RECT  5.17 4.735 8.515 4.74 ;
      RECT  5.165 4.74 8.515 4.745 ;
      RECT  5.16 4.745 8.515 4.75 ;
      RECT  5.155 4.75 8.515 4.755 ;
      RECT  5.15 4.755 8.515 4.76 ;
      RECT  5.145 4.76 8.515 4.765 ;
      RECT  5.14 4.765 8.515 4.77 ;
      RECT  5.135 4.77 8.515 4.775 ;
      RECT  5.13 4.775 8.515 4.78 ;
      RECT  5.125 4.78 8.515 4.785 ;
      RECT  5.12 4.785 8.515 4.79 ;
      RECT  5.115 4.79 8.515 4.795 ;
      RECT  5.11 4.795 8.515 4.8 ;
      RECT  5.105 4.8 8.515 4.805 ;
      RECT  5.1 4.805 8.515 4.81 ;
      RECT  5.095 4.81 8.515 4.815 ;
      RECT  5.09 4.815 8.515 4.82 ;
      RECT  5.085 4.82 8.515 4.825 ;
      RECT  5.08 4.825 8.515 4.83 ;
      RECT  5.075 4.83 8.515 4.835 ;
      RECT  5.07 4.835 8.515 4.84 ;
      RECT  5.065 4.84 8.515 4.845 ;
      RECT  5.06 4.845 8.515 4.85 ;
      RECT  5.055 4.85 8.515 4.855 ;
      RECT  5.05 4.855 8.515 4.86 ;
      RECT  5.045 4.86 8.515 4.865 ;
      RECT  5.04 4.865 8.515 4.87 ;
      RECT  5.035 4.87 8.515 4.875 ;
      RECT  5.03 4.875 8.515 4.88 ;
      RECT  5.025 4.88 8.515 4.885 ;
      RECT  5.02 4.885 8.515 4.89 ;
      RECT  5.015 4.89 8.515 4.895 ;
      RECT  5.01 4.895 5.335 4.9 ;
      RECT  8.285 4.895 8.515 5.0 ;
      RECT  5.005 4.9 5.33 4.905 ;
      RECT  5.0 4.905 5.325 4.91 ;
      RECT  4.995 4.91 5.32 4.915 ;
      RECT  4.99 4.915 5.315 4.92 ;
      RECT  4.985 4.92 5.31 4.925 ;
      RECT  4.98 4.925 5.305 4.93 ;
      RECT  4.975 4.93 5.3 4.935 ;
      RECT  4.97 4.935 5.295 4.94 ;
      RECT  4.965 4.94 5.29 4.945 ;
      RECT  4.96 4.945 5.285 4.95 ;
      RECT  4.955 4.95 5.28 4.955 ;
      RECT  4.95 4.955 5.275 4.96 ;
      RECT  4.945 4.96 5.27 4.965 ;
      RECT  4.94 4.965 5.265 4.97 ;
      RECT  4.935 4.97 5.26 4.975 ;
      RECT  4.93 4.975 5.255 4.98 ;
      RECT  4.925 4.98 5.25 4.985 ;
      RECT  4.92 4.985 5.245 4.99 ;
      RECT  4.915 4.99 5.24 4.995 ;
      RECT  4.91 4.995 5.235 5.0 ;
      RECT  0.18 4.365 1.74 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 5.23 5.005 ;
      RECT  8.285 5.0 10.81 5.23 ;
      RECT  1.51 5.005 5.225 5.01 ;
      RECT  1.51 5.01 5.22 5.015 ;
      RECT  1.51 5.015 5.215 5.02 ;
      RECT  1.51 5.02 5.21 5.025 ;
      RECT  1.51 5.025 5.205 5.03 ;
      RECT  1.51 5.03 5.2 5.035 ;
      RECT  1.51 5.035 5.195 5.04 ;
      RECT  1.51 5.04 5.19 5.045 ;
      RECT  1.51 5.045 5.185 5.05 ;
      RECT  1.51 5.05 5.18 5.055 ;
      RECT  1.51 5.055 5.175 5.06 ;
      RECT  1.51 5.06 5.17 5.065 ;
      RECT  1.51 5.065 5.165 5.07 ;
      RECT  1.51 5.07 5.16 5.075 ;
      RECT  1.51 5.075 5.155 5.08 ;
      RECT  1.51 5.08 5.15 5.085 ;
      RECT  1.51 5.085 5.145 5.09 ;
      RECT  1.51 5.09 5.14 5.095 ;
      RECT  1.51 5.095 5.135 5.1 ;
      RECT  1.51 5.1 5.13 5.105 ;
      RECT  1.51 5.105 5.125 5.11 ;
      RECT  1.51 5.11 5.12 5.115 ;
      RECT  1.51 5.115 5.115 5.12 ;
      RECT  1.51 5.12 5.11 5.125 ;
      RECT  1.51 5.125 5.105 5.13 ;
      RECT  1.51 5.13 5.1 5.135 ;
      RECT  1.51 5.135 5.095 5.14 ;
      RECT  1.51 5.14 5.09 5.145 ;
      RECT  1.51 5.145 5.085 5.15 ;
      RECT  1.51 5.15 5.08 5.155 ;
      RECT  1.51 5.155 5.075 5.16 ;
      RECT  1.51 5.16 5.07 5.165 ;
      RECT  1.51 5.165 5.065 5.17 ;
      RECT  1.51 5.17 5.06 5.175 ;
      RECT  1.51 5.175 5.055 5.18 ;
      RECT  1.51 5.18 5.05 5.185 ;
      RECT  1.51 5.185 5.045 5.19 ;
      RECT  1.51 5.19 5.04 5.195 ;
      RECT  1.51 5.195 5.035 5.2 ;
      RECT  1.51 5.2 5.03 5.205 ;
      RECT  1.51 5.205 5.025 5.21 ;
      RECT  1.51 5.21 5.02 5.215 ;
      RECT  1.51 5.215 5.015 5.22 ;
      RECT  1.51 5.22 5.01 5.225 ;
      RECT  1.51 5.225 5.005 5.23 ;
  END
END MDN_FDNSBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FDP_4
#      Description : D-Flip Flop, pos-edge triggered
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDP_4
  CLASS CORE ;
  FOREIGN MDN_FDP_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 4.365 0.7 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.92 1.565 16.2 1.795 ;
      RECT  15.565 1.795 15.795 3.245 ;
      RECT  12.92 3.245 16.2 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.1 1.565 22.22 1.795 ;
      RECT  20.045 1.795 20.275 3.245 ;
      RECT  18.1 3.245 22.22 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.03 5.46 12.435 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.925 -0.14 19.6 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  14.445 -0.14 16.915 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  11.03 -0.14 12.435 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  2.8 -0.14 3.92 0.14 ;
      RECT  3.19 0.14 3.53 0.465 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.485 0.37 7.45 0.6 ;
      RECT  5.485 0.6 5.715 0.73 ;
      RECT  8.23 0.37 11.61 0.6 ;
      RECT  11.38 0.6 11.61 1.005 ;
      RECT  11.38 1.005 12.435 1.235 ;
      RECT  12.205 1.235 12.435 2.415 ;
      RECT  12.205 2.415 15.29 2.645 ;
      RECT  12.205 2.645 12.435 4.365 ;
      RECT  11.38 4.365 12.435 4.595 ;
      RECT  17.19 0.37 17.53 0.6 ;
      RECT  17.19 0.6 17.42 1.005 ;
      RECT  14.95 0.37 16.415 0.6 ;
      RECT  16.185 0.6 16.415 1.005 ;
      RECT  16.185 1.005 17.42 1.235 ;
      RECT  19.43 0.37 20.89 0.6 ;
      RECT  2.62 0.37 2.96 0.715 ;
      RECT  1.465 0.715 5.21 0.945 ;
      RECT  4.87 0.37 5.21 0.715 ;
      RECT  1.465 0.945 1.695 1.005 ;
      RECT  0.18 1.005 1.695 1.235 ;
      RECT  0.445 1.235 0.675 3.245 ;
      RECT  0.18 3.245 0.675 3.475 ;
      RECT  5.485 1.005 6.54 1.235 ;
      RECT  5.485 1.235 5.715 1.74 ;
      RECT  3.96 1.74 5.715 1.97 ;
      RECT  8.44 1.005 11.02 1.235 ;
      RECT  1.96 1.22 5.0 1.45 ;
      RECT  1.96 1.45 2.19 1.565 ;
      RECT  1.72 1.565 2.19 1.795 ;
      RECT  6.9 1.465 9.635 1.695 ;
      RECT  9.405 1.695 9.635 1.975 ;
      RECT  9.405 1.975 10.195 2.205 ;
      RECT  9.965 2.205 10.195 3.245 ;
      RECT  7.725 3.245 11.02 3.475 ;
      RECT  7.725 3.475 7.955 3.805 ;
      RECT  6.8 3.805 7.955 4.035 ;
      RECT  6.8 4.035 7.03 4.365 ;
      RECT  4.365 4.365 7.03 4.595 ;
      RECT  4.365 4.595 4.595 5.0 ;
      RECT  3.75 5.0 4.595 5.23 ;
      RECT  9.91 1.5 11.875 1.73 ;
      RECT  11.645 1.73 11.875 3.805 ;
      RECT  9.91 3.805 11.875 4.035 ;
      RECT  17.245 1.565 17.74 1.795 ;
      RECT  17.245 1.795 17.475 2.685 ;
      RECT  17.245 2.685 19.715 2.915 ;
      RECT  18.365 2.36 18.595 2.685 ;
      RECT  19.485 2.36 19.715 2.685 ;
      RECT  17.245 2.915 17.475 3.245 ;
      RECT  17.245 3.245 17.74 3.475 ;
      RECT  6.045 1.93 8.515 2.16 ;
      RECT  8.285 2.16 8.515 2.44 ;
      RECT  6.045 2.16 6.275 2.685 ;
      RECT  8.285 2.44 9.69 2.67 ;
      RECT  2.42 1.68 3.475 1.91 ;
      RECT  3.245 1.91 3.475 2.685 ;
      RECT  3.245 2.685 6.275 2.915 ;
      RECT  3.245 2.915 3.475 3.805 ;
      RECT  2.42 3.805 3.475 4.035 ;
      RECT  20.605 2.36 20.835 2.685 ;
      RECT  20.605 2.685 21.955 2.915 ;
      RECT  21.725 2.36 21.955 2.685 ;
      RECT  7.165 2.39 7.395 3.245 ;
      RECT  5.43 3.245 7.395 3.475 ;
      RECT  3.96 3.245 5.0 3.475 ;
      RECT  3.805 3.805 6.54 4.035 ;
      RECT  3.805 4.035 4.035 4.365 ;
      RECT  1.72 4.365 4.035 4.595 ;
      RECT  8.44 3.805 9.48 4.035 ;
      RECT  7.26 4.365 10.195 4.595 ;
      RECT  7.26 4.595 7.49 5.0 ;
      RECT  9.965 4.595 10.195 5.0 ;
      RECT  4.87 5.0 7.49 5.23 ;
      RECT  9.965 5.0 10.81 5.23 ;
  END
END MDN_FDP_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FDP_1
#      Description : D-Flip Flop, pos-edge triggered
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDP_1
  CLASS CORE ;
  FOREIGN MDN_FDP_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 4.365 0.7 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.62 1.005 14.115 1.235 ;
      RECT  13.885 1.235 14.115 3.245 ;
      RECT  13.62 3.245 14.115 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.765 1.565 13.26 1.795 ;
      RECT  12.765 1.795 12.995 3.805 ;
      RECT  12.765 3.805 13.26 4.035 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.935 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  6.55 5.46 7.955 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  2.8 -0.14 3.92 0.14 ;
      RECT  3.19 0.14 3.53 0.465 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.37 7.45 0.6 ;
      RECT  12.765 0.37 14.17 0.6 ;
      RECT  12.765 0.6 12.995 1.005 ;
      RECT  8.23 0.37 11.665 0.6 ;
      RECT  11.435 0.6 11.665 1.005 ;
      RECT  11.435 1.005 12.995 1.235 ;
      RECT  12.205 1.235 12.435 4.015 ;
      RECT  11.38 4.015 12.435 4.245 ;
      RECT  1.775 0.695 4.945 0.925 ;
      RECT  1.775 0.925 2.005 1.29 ;
      RECT  4.715 0.925 4.945 1.29 ;
      RECT  8.44 1.005 11.02 1.235 ;
      RECT  2.42 1.155 3.475 1.385 ;
      RECT  3.245 1.385 3.475 1.985 ;
      RECT  3.245 1.985 8.515 2.215 ;
      RECT  8.285 2.215 8.515 2.445 ;
      RECT  6.045 2.215 6.275 2.995 ;
      RECT  8.285 2.445 9.465 2.675 ;
      RECT  3.245 2.995 6.275 3.225 ;
      RECT  3.245 3.225 3.475 3.805 ;
      RECT  2.42 3.805 3.475 4.035 ;
      RECT  9.96 1.51 11.875 1.74 ;
      RECT  11.645 1.74 11.875 3.555 ;
      RECT  9.91 3.555 11.875 3.785 ;
      RECT  10.525 3.785 10.755 4.475 ;
      RECT  10.525 4.475 12.94 4.705 ;
      RECT  12.71 4.705 12.94 5.0 ;
      RECT  11.59 4.705 11.93 5.23 ;
      RECT  12.71 5.0 13.05 5.23 ;
      RECT  3.96 1.525 6.54 1.755 ;
      RECT  6.9 1.525 9.635 1.755 ;
      RECT  9.405 1.755 9.635 1.985 ;
      RECT  9.405 1.985 10.195 2.215 ;
      RECT  9.965 2.215 10.195 3.095 ;
      RECT  7.725 3.095 11.02 3.325 ;
      RECT  7.725 3.325 7.955 3.925 ;
      RECT  6.795 3.925 7.955 4.155 ;
      RECT  6.795 4.155 7.025 4.44 ;
      RECT  4.365 4.44 7.025 4.67 ;
      RECT  4.365 4.67 4.595 5.0 ;
      RECT  3.75 5.0 4.595 5.23 ;
      RECT  0.18 1.625 2.915 1.855 ;
      RECT  2.685 1.855 2.915 2.445 ;
      RECT  0.445 1.855 0.675 3.245 ;
      RECT  2.685 2.445 5.21 2.675 ;
      RECT  0.18 3.245 0.675 3.475 ;
      RECT  7.11 2.445 7.45 2.675 ;
      RECT  7.165 2.675 7.395 3.465 ;
      RECT  5.43 3.465 7.395 3.695 ;
      RECT  3.96 3.465 5.0 3.695 ;
      RECT  8.44 3.805 9.48 4.035 ;
      RECT  3.805 3.935 6.54 4.165 ;
      RECT  3.805 4.165 4.035 4.365 ;
      RECT  1.72 4.365 4.035 4.595 ;
      RECT  7.255 4.39 10.195 4.62 ;
      RECT  7.255 4.62 7.485 5.0 ;
      RECT  9.965 4.62 10.195 5.0 ;
      RECT  4.87 5.0 7.485 5.23 ;
      RECT  9.965 5.0 10.81 5.23 ;
  END
END MDN_FDP_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FDP_2
#      Description : D-Flip Flop, pos-edge triggered
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDP_2
  CLASS CORE ;
  FOREIGN MDN_FDP_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 4.365 0.7 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.16 1.565 16.2 1.795 ;
      RECT  15.565 1.795 15.795 3.245 ;
      RECT  15.16 3.245 16.2 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.92 1.565 13.96 1.795 ;
      RECT  13.325 1.795 13.555 3.245 ;
      RECT  12.92 3.245 13.96 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  12.205 4.94 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  6.55 5.46 7.955 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  11.76 -0.14 12.435 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  2.8 -0.14 3.92 0.14 ;
      RECT  3.19 0.14 3.53 0.475 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.37 7.45 0.6 ;
      RECT  14.95 0.37 16.41 0.6 ;
      RECT  15.005 0.6 15.235 1.005 ;
      RECT  8.225 0.37 11.61 0.6 ;
      RECT  11.38 0.6 11.61 1.005 ;
      RECT  11.38 1.005 15.235 1.235 ;
      RECT  12.205 1.235 12.435 4.02 ;
      RECT  11.38 4.02 12.435 4.25 ;
      RECT  1.775 0.705 4.945 0.935 ;
      RECT  1.775 0.935 2.005 1.29 ;
      RECT  4.715 0.935 4.945 1.29 ;
      RECT  0.18 1.005 0.675 1.235 ;
      RECT  0.445 1.235 0.675 1.63 ;
      RECT  0.445 1.63 2.915 1.86 ;
      RECT  2.685 1.86 2.915 2.44 ;
      RECT  0.445 1.86 0.675 3.245 ;
      RECT  2.685 2.44 5.215 2.67 ;
      RECT  0.18 3.245 0.675 3.475 ;
      RECT  8.44 1.005 11.02 1.235 ;
      RECT  2.42 1.17 3.475 1.4 ;
      RECT  3.245 1.4 3.475 1.98 ;
      RECT  3.245 1.98 8.515 2.21 ;
      RECT  8.285 2.21 8.515 2.445 ;
      RECT  6.045 2.21 6.275 2.9 ;
      RECT  8.285 2.445 9.69 2.675 ;
      RECT  3.245 2.9 6.275 3.13 ;
      RECT  3.245 3.13 3.475 3.805 ;
      RECT  2.42 3.805 3.475 4.035 ;
      RECT  9.91 1.49 11.875 1.72 ;
      RECT  11.645 1.72 11.875 3.56 ;
      RECT  9.86 3.56 11.875 3.79 ;
      RECT  10.525 3.79 10.755 4.48 ;
      RECT  10.525 4.48 12.94 4.71 ;
      RECT  12.71 4.71 12.94 5.0 ;
      RECT  11.59 4.71 11.93 5.23 ;
      RECT  12.71 5.0 14.17 5.23 ;
      RECT  6.9 1.51 9.425 1.74 ;
      RECT  9.195 1.74 9.425 1.965 ;
      RECT  9.195 1.965 10.195 2.195 ;
      RECT  9.965 2.195 10.195 3.095 ;
      RECT  7.725 3.095 11.02 3.325 ;
      RECT  7.725 3.325 7.955 3.82 ;
      RECT  6.775 3.82 7.955 4.05 ;
      RECT  6.775 4.05 7.005 4.44 ;
      RECT  4.365 4.44 7.005 4.67 ;
      RECT  4.365 4.67 4.595 5.0 ;
      RECT  3.75 5.0 4.595 5.23 ;
      RECT  3.96 1.52 6.54 1.75 ;
      RECT  6.605 2.44 7.45 2.67 ;
      RECT  6.605 2.67 6.835 3.36 ;
      RECT  5.43 3.36 6.835 3.59 ;
      RECT  3.96 3.465 5.0 3.695 ;
      RECT  8.44 3.805 9.48 4.035 ;
      RECT  3.805 3.935 6.54 4.165 ;
      RECT  3.805 4.165 4.035 4.365 ;
      RECT  1.72 4.365 4.035 4.595 ;
      RECT  7.255 4.365 10.195 4.595 ;
      RECT  7.255 4.595 7.485 5.0 ;
      RECT  9.965 4.595 10.195 5.0 ;
      RECT  4.87 5.0 7.485 5.23 ;
      RECT  9.965 5.0 10.81 5.23 ;
  END
END MDN_FDP_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPHRBQ_1
#      Description : D-Flip Flop, pos-edge triggered, lo-async-clear, sync hold, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D&!EN)|(iq&EN),clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPHRBQ_1
  CLASS CORE ;
  FOREIGN MDN_FDPHRBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 4.365 6.3 5.0 ;
      RECT  5.99 5.0 6.33 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.485 1.565 19.98 1.795 ;
      RECT  19.485 1.795 19.715 3.245 ;
      RECT  19.485 3.245 19.98 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.22 2.125 17.5 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.87 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.99 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  -0.17 5.46 0.56 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  17.245 -0.14 17.92 0.14 ;
      RECT  17.245 0.14 17.475 1.005 ;
      RECT  17.245 1.005 17.74 1.235 ;
      RECT  12.765 -0.14 14.0 0.14 ;
      RECT  12.765 0.14 12.995 1.005 ;
      RECT  12.765 1.005 13.26 1.235 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  1.68 -0.14 2.8 0.14 ;
      RECT  2.125 0.14 2.355 1.005 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  2.63 0.37 3.475 0.6 ;
      RECT  3.245 0.6 3.475 0.98 ;
      RECT  3.17 0.98 3.55 1.26 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  8.23 0.37 10.25 0.6 ;
      RECT  11.59 0.37 11.93 0.6 ;
      RECT  11.7 0.6 11.93 1.005 ;
      RECT  9.965 1.005 12.435 1.235 ;
      RECT  9.965 1.235 10.195 1.465 ;
      RECT  12.205 1.235 12.435 1.525 ;
      RECT  7.99 1.465 10.195 1.695 ;
      RECT  12.205 1.525 15.5 1.755 ;
      RECT  7.99 1.695 8.22 3.03 ;
      RECT  15.27 1.755 15.5 3.08 ;
      RECT  7.99 3.03 8.78 3.26 ;
      RECT  15.16 3.08 15.5 3.31 ;
      RECT  14.39 0.37 16.41 0.6 ;
      RECT  13.49 0.98 13.87 1.005 ;
      RECT  13.49 1.005 16.915 1.235 ;
      RECT  13.49 1.235 13.87 1.26 ;
      RECT  16.685 1.235 16.915 1.565 ;
      RECT  16.685 1.565 18.44 1.795 ;
      RECT  16.685 1.795 16.915 3.54 ;
      RECT  13.62 3.54 18.44 3.77 ;
      RECT  3.805 1.005 9.48 1.235 ;
      RECT  3.805 1.235 4.035 1.565 ;
      RECT  5.485 1.235 5.715 3.81 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 1.565 ;
      RECT  1.005 1.565 4.035 1.795 ;
      RECT  1.005 1.795 1.235 3.53 ;
      RECT  5.485 3.81 6.835 3.95 ;
      RECT  5.485 3.95 11.02 4.04 ;
      RECT  6.605 4.04 11.02 4.18 ;
      RECT  10.68 1.47 11.72 1.7 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 3.245 ;
      RECT  1.565 2.35 1.795 2.685 ;
      RECT  1.565 2.685 3.475 2.915 ;
      RECT  3.245 2.915 3.475 3.245 ;
      RECT  3.245 3.245 5.155 3.475 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 2.685 ;
      RECT  6.045 2.685 7.3 2.915 ;
      RECT  7.07 2.39 7.3 2.685 ;
      RECT  6.045 2.915 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
      RECT  15.86 1.565 16.355 1.795 ;
      RECT  16.125 1.795 16.355 3.08 ;
      RECT  15.86 3.08 16.355 3.31 ;
      RECT  9.47 1.985 15.025 2.215 ;
      RECT  14.795 2.215 15.025 2.655 ;
      RECT  9.47 2.215 9.7 2.69 ;
      RECT  8.45 2.405 9.24 2.635 ;
      RECT  9.01 2.635 9.24 3.03 ;
      RECT  9.01 3.03 10.25 3.26 ;
      RECT  10.47 2.445 14.17 2.675 ;
      RECT  10.525 2.675 10.755 3.49 ;
      RECT  6.9 1.565 7.76 1.795 ;
      RECT  7.53 1.795 7.76 3.245 ;
      RECT  6.9 3.245 7.76 3.475 ;
      RECT  7.53 3.475 7.76 3.49 ;
      RECT  7.53 3.49 10.755 3.72 ;
      RECT  1.72 3.245 2.76 3.475 ;
      RECT  15.86 4.07 18.035 4.3 ;
      RECT  17.805 4.3 18.035 4.365 ;
      RECT  17.805 4.365 19.66 4.595 ;
      RECT  18.42 4.595 18.65 5.0 ;
      RECT  19.43 4.595 19.66 5.0 ;
      RECT  18.31 5.0 18.65 5.23 ;
      RECT  19.43 5.0 19.77 5.23 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  7.22 4.41 8.515 4.64 ;
      RECT  7.22 4.64 7.45 5.0 ;
      RECT  8.285 4.64 8.515 5.0 ;
      RECT  7.11 5.0 7.45 5.23 ;
      RECT  8.285 5.0 9.69 5.23 ;
      RECT  9.14 4.41 13.26 4.64 ;
      RECT  13.885 4.53 17.42 4.76 ;
      RECT  13.885 4.76 14.115 5.0 ;
      RECT  17.19 4.76 17.42 5.0 ;
      RECT  12.71 5.0 14.115 5.23 ;
      RECT  17.19 5.0 17.53 5.23 ;
      RECT  14.39 5.0 16.41 5.23 ;
      LAYER METAL2 ;
      RECT  3.17 0.98 13.87 1.26 ;
      LAYER VIA12 ;
      RECT  3.23 0.99 3.49 1.25 ;
      RECT  13.55 0.99 13.81 1.25 ;
  END
END MDN_FDPHRBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPHRBQ_2
#      Description : D-Flip Flop, pos-edge triggered, lo-async-clear, sync hold, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D&!EN)|(iq&EN),clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPHRBQ_2
  CLASS CORE ;
  FOREIGN MDN_FDPHRBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 4.365 6.3 5.0 ;
      RECT  5.99 5.0 6.33 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.64 1.565 20.68 1.795 ;
      RECT  20.045 1.795 20.275 3.245 ;
      RECT  19.64 3.245 20.68 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.22 2.125 17.5 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.87 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.92 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  12.205 4.875 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  -0.17 5.46 0.56 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.8 -0.14 17.475 0.14 ;
      RECT  17.245 0.14 17.475 1.005 ;
      RECT  17.245 1.005 17.74 1.235 ;
      RECT  12.765 -0.14 14.0 0.14 ;
      RECT  12.765 0.14 12.995 1.005 ;
      RECT  12.765 1.005 13.26 1.235 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  1.68 -0.14 2.8 0.14 ;
      RECT  2.125 0.14 2.355 1.0 ;
      RECT  1.72 1.0 2.76 1.23 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  2.63 0.37 3.475 0.6 ;
      RECT  3.245 0.6 3.475 0.98 ;
      RECT  3.17 0.98 3.55 1.26 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  8.23 0.37 10.25 0.6 ;
      RECT  11.59 0.37 11.93 0.6 ;
      RECT  11.59 0.6 11.82 1.005 ;
      RECT  9.965 1.005 12.435 1.235 ;
      RECT  9.965 1.235 10.195 1.47 ;
      RECT  12.205 1.235 12.435 1.49 ;
      RECT  7.915 1.47 10.195 1.7 ;
      RECT  12.205 1.49 15.53 1.72 ;
      RECT  7.915 1.7 8.145 3.03 ;
      RECT  15.3 1.72 15.53 3.07 ;
      RECT  7.915 3.03 8.78 3.26 ;
      RECT  15.16 3.07 15.53 3.3 ;
      RECT  14.39 0.37 16.41 0.6 ;
      RECT  13.49 0.98 13.87 1.005 ;
      RECT  13.49 1.005 16.915 1.235 ;
      RECT  13.49 1.235 13.87 1.26 ;
      RECT  16.685 1.235 16.915 1.565 ;
      RECT  16.685 1.565 18.44 1.795 ;
      RECT  16.685 1.795 16.915 3.245 ;
      RECT  16.685 3.245 18.44 3.475 ;
      RECT  16.685 3.475 16.915 3.535 ;
      RECT  15.005 3.535 16.915 3.765 ;
      RECT  15.005 3.765 15.235 3.805 ;
      RECT  13.62 3.805 15.235 4.035 ;
      RECT  3.8 1.005 9.48 1.235 ;
      RECT  3.8 1.235 4.03 1.565 ;
      RECT  5.485 1.235 5.715 3.805 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 1.565 ;
      RECT  1.005 1.565 4.03 1.795 ;
      RECT  1.005 1.795 1.235 3.53 ;
      RECT  5.485 3.805 7.19 3.95 ;
      RECT  5.485 3.95 11.02 4.035 ;
      RECT  6.96 4.035 11.02 4.18 ;
      RECT  10.68 1.47 11.72 1.7 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 3.245 ;
      RECT  1.565 2.35 1.795 2.685 ;
      RECT  1.565 2.685 3.475 2.915 ;
      RECT  3.245 2.915 3.475 3.245 ;
      RECT  3.245 3.245 5.155 3.475 ;
      RECT  15.86 1.565 16.355 1.795 ;
      RECT  16.125 1.795 16.355 3.075 ;
      RECT  15.86 3.075 16.355 3.305 ;
      RECT  9.47 1.95 15.065 2.18 ;
      RECT  9.47 2.18 9.7 2.69 ;
      RECT  14.835 2.18 15.065 2.69 ;
      RECT  6.255 1.51 6.485 2.405 ;
      RECT  6.255 2.405 7.225 2.635 ;
      RECT  6.255 2.635 6.485 3.53 ;
      RECT  8.375 2.405 9.24 2.635 ;
      RECT  9.01 2.635 9.24 3.03 ;
      RECT  9.01 3.03 10.25 3.26 ;
      RECT  10.47 2.445 14.17 2.675 ;
      RECT  10.525 2.675 10.755 3.49 ;
      RECT  6.9 1.565 7.685 1.795 ;
      RECT  7.455 1.795 7.685 3.245 ;
      RECT  6.9 3.245 7.685 3.475 ;
      RECT  7.455 3.475 7.685 3.49 ;
      RECT  7.455 3.49 10.755 3.72 ;
      RECT  1.72 3.245 2.76 3.475 ;
      RECT  15.86 4.0 18.035 4.23 ;
      RECT  17.805 4.23 18.035 4.365 ;
      RECT  17.805 4.365 19.66 4.595 ;
      RECT  18.42 4.595 18.65 5.0 ;
      RECT  19.43 4.595 19.66 5.0 ;
      RECT  18.31 5.0 18.65 5.23 ;
      RECT  19.43 5.0 20.89 5.23 ;
      RECT  2.685 4.365 4.3 4.595 ;
      RECT  2.685 4.595 2.915 4.925 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 4.925 ;
      RECT  0.445 4.925 2.915 5.155 ;
      RECT  7.22 4.41 8.515 4.64 ;
      RECT  7.22 4.64 7.45 5.0 ;
      RECT  8.285 4.64 8.515 5.0 ;
      RECT  7.11 5.0 7.45 5.23 ;
      RECT  8.285 5.0 9.69 5.23 ;
      RECT  9.14 4.415 13.26 4.645 ;
      RECT  13.885 4.46 17.42 4.69 ;
      RECT  13.885 4.69 14.115 5.0 ;
      RECT  17.19 4.69 17.42 5.0 ;
      RECT  12.71 5.0 14.115 5.23 ;
      RECT  17.19 5.0 17.53 5.23 ;
      RECT  14.39 5.0 16.41 5.23 ;
      LAYER METAL2 ;
      RECT  3.17 0.98 13.87 1.26 ;
      LAYER VIA12 ;
      RECT  3.23 0.99 3.49 1.25 ;
      RECT  13.55 0.99 13.81 1.25 ;
  END
END MDN_FDPHRBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPHRBQ_4
#      Description : D-Flip Flop, pos-edge triggered, lo-async-clear, sync hold, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D&!EN)|(iq&EN),clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPHRBQ_4
  CLASS CORE ;
  FOREIGN MDN_FDPHRBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 24.64 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 4.365 6.3 5.0 ;
      RECT  5.99 5.0 6.33 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.64 1.565 22.92 1.795 ;
      RECT  20.045 1.795 20.275 3.245 ;
      RECT  19.64 3.245 22.925 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.22 2.125 17.5 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.81 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  20.72 5.46 21.395 5.74 ;
      RECT  18.925 4.87 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.99 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  -0.17 5.46 0.56 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 24.64 5.74 ;
      LAYER VIA12 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  24.23 5.47 24.49 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 -0.14 24.81 0.14 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  20.72 -0.14 21.395 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.8 -0.14 17.475 0.14 ;
      RECT  17.245 0.14 17.475 1.005 ;
      RECT  17.245 1.005 17.74 1.235 ;
      RECT  12.765 -0.14 14.0 0.14 ;
      RECT  12.765 0.14 12.995 1.005 ;
      RECT  12.765 1.005 13.26 1.235 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  1.68 -0.14 2.8 0.14 ;
      RECT  2.125 0.14 2.355 1.005 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 24.64 0.14 ;
      LAYER VIA12 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  20.87 -0.13 21.13 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 8.57 0.445 ;
      RECT  8.23 0.445 10.25 0.675 ;
      RECT  16.07 0.37 16.41 0.445 ;
      RECT  14.39 0.445 16.41 0.675 ;
      RECT  2.63 0.37 3.475 0.6 ;
      RECT  3.245 0.6 3.475 0.98 ;
      RECT  3.17 0.98 3.55 1.26 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  11.59 0.37 11.93 0.6 ;
      RECT  11.59 0.6 11.82 0.95 ;
      RECT  9.965 0.95 12.435 1.18 ;
      RECT  9.965 1.18 10.195 1.465 ;
      RECT  12.205 1.18 12.435 1.49 ;
      RECT  7.995 1.465 10.195 1.695 ;
      RECT  12.205 1.49 15.63 1.72 ;
      RECT  7.995 1.695 8.225 3.03 ;
      RECT  15.4 1.72 15.63 3.075 ;
      RECT  7.995 3.03 8.78 3.26 ;
      RECT  15.16 3.075 15.63 3.305 ;
      RECT  13.49 0.98 13.87 1.005 ;
      RECT  13.49 1.005 16.915 1.235 ;
      RECT  13.49 1.235 13.87 1.26 ;
      RECT  16.685 1.235 16.915 1.565 ;
      RECT  16.685 1.565 18.44 1.795 ;
      RECT  16.685 1.795 16.915 3.535 ;
      RECT  13.62 3.535 18.44 3.765 ;
      RECT  3.805 1.005 9.48 1.235 ;
      RECT  3.805 1.235 4.035 1.565 ;
      RECT  5.485 1.235 5.715 3.805 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 1.565 ;
      RECT  1.005 1.565 4.035 1.795 ;
      RECT  1.005 1.795 1.235 3.53 ;
      RECT  5.485 3.805 6.835 3.95 ;
      RECT  5.485 3.95 11.02 4.035 ;
      RECT  6.605 4.035 11.02 4.18 ;
      RECT  10.68 1.46 11.72 1.69 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 3.245 ;
      RECT  1.565 2.35 1.795 2.685 ;
      RECT  1.565 2.685 3.475 2.915 ;
      RECT  3.245 2.915 3.475 3.245 ;
      RECT  3.245 3.245 5.155 3.475 ;
      RECT  15.86 1.565 16.355 1.795 ;
      RECT  16.125 1.795 16.355 3.075 ;
      RECT  15.86 3.075 16.355 3.305 ;
      RECT  9.47 1.95 15.165 2.18 ;
      RECT  9.47 2.18 9.7 2.69 ;
      RECT  14.935 2.18 15.165 2.69 ;
      RECT  6.255 1.51 6.485 2.4 ;
      RECT  6.255 2.4 7.26 2.63 ;
      RECT  6.255 2.63 6.485 3.53 ;
      RECT  8.455 2.405 9.24 2.635 ;
      RECT  9.01 2.635 9.24 3.03 ;
      RECT  9.01 3.03 10.2 3.26 ;
      RECT  10.47 2.445 14.17 2.675 ;
      RECT  10.525 2.675 10.755 3.49 ;
      RECT  6.9 1.565 7.765 1.795 ;
      RECT  7.535 1.795 7.765 3.245 ;
      RECT  6.9 3.245 7.765 3.475 ;
      RECT  7.535 3.475 7.765 3.49 ;
      RECT  7.535 3.49 10.755 3.72 ;
      RECT  20.605 2.35 20.835 2.685 ;
      RECT  20.605 2.685 23.075 2.915 ;
      RECT  21.725 2.35 21.955 2.685 ;
      RECT  22.845 2.35 23.075 2.685 ;
      RECT  1.72 3.245 2.76 3.475 ;
      RECT  15.86 4.07 18.035 4.3 ;
      RECT  17.805 4.3 18.035 4.365 ;
      RECT  17.805 4.365 19.66 4.595 ;
      RECT  18.42 4.595 18.65 5.0 ;
      RECT  19.43 4.595 19.66 5.0 ;
      RECT  18.31 5.0 18.65 5.23 ;
      RECT  19.43 5.0 20.89 5.23 ;
      RECT  2.685 4.365 4.3 4.595 ;
      RECT  2.685 4.595 2.915 4.925 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 4.925 ;
      RECT  0.445 4.925 2.915 5.155 ;
      RECT  7.22 4.41 8.515 4.64 ;
      RECT  7.22 4.64 7.45 5.0 ;
      RECT  8.285 4.64 8.515 5.0 ;
      RECT  7.11 5.0 7.45 5.23 ;
      RECT  8.285 5.0 9.69 5.23 ;
      RECT  9.14 4.41 13.26 4.64 ;
      RECT  13.885 4.53 17.42 4.76 ;
      RECT  13.885 4.76 14.115 5.0 ;
      RECT  17.19 4.76 17.42 5.0 ;
      RECT  12.71 5.0 14.115 5.23 ;
      RECT  17.19 5.0 17.53 5.23 ;
      RECT  14.39 5.0 16.41 5.23 ;
      LAYER METAL2 ;
      RECT  3.17 0.98 13.87 1.26 ;
      LAYER VIA12 ;
      RECT  3.23 0.99 3.49 1.25 ;
      RECT  13.55 0.99 13.81 1.25 ;
  END
END MDN_FDPHRBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPQ_1
#      Description : D-Flip Flop, pos-edge triggered, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPQ_1
  CLASS CORE ;
  FOREIGN MDN_FDPQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 4.365 11.9 5.0 ;
      RECT  11.59 5.0 11.93 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.765 1.565 13.26 1.795 ;
      RECT  12.765 1.795 12.995 3.245 ;
      RECT  12.765 3.245 13.26 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  5.485 5.08 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.66 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  5.48 1.005 6.22 1.235 ;
      RECT  5.48 1.235 5.71 1.565 ;
      RECT  3.19 1.565 5.715 1.795 ;
      RECT  4.365 1.795 4.595 3.03 ;
      RECT  3.19 3.03 4.595 3.26 ;
      RECT  10.47 0.37 10.81 0.6 ;
      RECT  10.47 0.6 10.7 1.005 ;
      RECT  7.725 1.005 10.7 1.235 ;
      RECT  7.725 1.235 7.955 3.315 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  10.93 1.005 12.94 1.235 ;
      RECT  10.93 1.235 11.16 1.51 ;
      RECT  10.735 1.51 11.16 1.795 ;
      RECT  10.735 1.795 10.965 2.405 ;
      RECT  9.35 2.405 10.965 2.635 ;
      RECT  10.735 2.635 10.965 3.46 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.005 5.0 1.235 ;
      RECT  1.72 1.565 2.835 1.57 ;
      RECT  1.72 1.57 2.915 1.795 ;
      RECT  2.685 1.795 2.915 2.415 ;
      RECT  2.685 2.415 4.09 2.645 ;
      RECT  2.685 2.645 2.915 3.03 ;
      RECT  1.72 3.03 2.915 3.26 ;
      RECT  6.045 1.565 7.24 1.795 ;
      RECT  6.045 1.795 6.275 2.405 ;
      RECT  4.87 2.405 6.275 2.635 ;
      RECT  6.045 2.635 6.275 3.7 ;
      RECT  6.045 3.7 7.095 3.93 ;
      RECT  6.865 3.93 7.095 4.01 ;
      RECT  6.865 4.01 8.78 4.24 ;
      RECT  8.44 1.565 9.48 1.795 ;
      RECT  11.435 1.51 11.875 1.85 ;
      RECT  11.645 1.85 11.875 3.805 ;
      RECT  9.405 3.805 11.875 4.035 ;
      RECT  9.405 4.035 9.635 4.54 ;
      RECT  4.565 4.16 6.635 4.39 ;
      RECT  4.565 4.39 4.795 4.54 ;
      RECT  6.405 4.39 6.635 4.54 ;
      RECT  2.74 4.54 4.795 4.77 ;
      RECT  6.405 4.54 9.635 4.77 ;
      RECT  2.74 4.77 2.97 5.0 ;
      RECT  8.23 4.77 8.46 5.0 ;
      RECT  1.51 5.0 2.97 5.23 ;
      RECT  8.23 5.0 8.57 5.23 ;
      RECT  8.285 3.245 9.48 3.475 ;
      RECT  8.285 3.475 8.515 3.545 ;
      RECT  6.895 3.235 7.32 3.24 ;
      RECT  6.895 3.24 7.325 3.245 ;
      RECT  6.895 3.245 7.33 3.25 ;
      RECT  6.895 3.25 7.335 3.255 ;
      RECT  6.895 3.255 7.34 3.26 ;
      RECT  6.895 3.26 7.345 3.265 ;
      RECT  6.895 3.265 7.35 3.27 ;
      RECT  6.895 3.27 7.355 3.275 ;
      RECT  6.895 3.275 7.36 3.28 ;
      RECT  6.895 3.28 7.365 3.285 ;
      RECT  6.895 3.285 7.37 3.29 ;
      RECT  6.895 3.29 7.375 3.295 ;
      RECT  6.895 3.295 7.38 3.3 ;
      RECT  6.895 3.3 7.385 3.305 ;
      RECT  6.895 3.305 7.39 3.31 ;
      RECT  6.895 3.31 7.395 3.315 ;
      RECT  6.895 3.315 7.4 3.32 ;
      RECT  6.895 3.32 7.405 3.325 ;
      RECT  6.895 3.325 7.41 3.33 ;
      RECT  6.895 3.33 7.415 3.335 ;
      RECT  6.895 3.335 7.42 3.34 ;
      RECT  6.895 3.34 7.425 3.345 ;
      RECT  6.895 3.345 7.43 3.35 ;
      RECT  6.895 3.35 7.435 3.355 ;
      RECT  6.895 3.355 7.44 3.36 ;
      RECT  6.895 3.36 7.445 3.365 ;
      RECT  6.895 3.365 7.45 3.37 ;
      RECT  6.895 3.37 7.455 3.375 ;
      RECT  6.895 3.375 7.46 3.38 ;
      RECT  6.895 3.38 7.465 3.385 ;
      RECT  6.895 3.385 7.47 3.39 ;
      RECT  6.895 3.39 7.475 3.395 ;
      RECT  6.895 3.395 7.48 3.4 ;
      RECT  6.895 3.4 7.485 3.405 ;
      RECT  6.895 3.405 7.49 3.41 ;
      RECT  6.895 3.41 7.495 3.415 ;
      RECT  6.895 3.415 7.5 3.42 ;
      RECT  6.895 3.42 7.505 3.425 ;
      RECT  6.895 3.425 7.51 3.43 ;
      RECT  6.895 3.43 7.515 3.435 ;
      RECT  6.895 3.435 7.52 3.44 ;
      RECT  6.895 3.44 7.525 3.445 ;
      RECT  6.895 3.445 7.53 3.45 ;
      RECT  6.895 3.45 7.535 3.455 ;
      RECT  6.895 3.455 7.54 3.46 ;
      RECT  6.895 3.46 7.545 3.465 ;
      RECT  7.215 3.465 7.55 3.47 ;
      RECT  7.22 3.47 7.555 3.475 ;
      RECT  7.225 3.475 7.56 3.48 ;
      RECT  7.23 3.48 7.565 3.485 ;
      RECT  7.235 3.485 7.57 3.49 ;
      RECT  7.24 3.49 7.575 3.495 ;
      RECT  7.245 3.495 7.58 3.5 ;
      RECT  7.25 3.5 7.585 3.505 ;
      RECT  7.255 3.505 7.59 3.51 ;
      RECT  7.26 3.51 7.595 3.515 ;
      RECT  7.265 3.515 7.6 3.52 ;
      RECT  7.27 3.52 7.605 3.525 ;
      RECT  7.275 3.525 7.61 3.53 ;
      RECT  7.28 3.53 7.615 3.535 ;
      RECT  7.285 3.535 7.62 3.54 ;
      RECT  7.29 3.54 7.625 3.545 ;
      RECT  7.295 3.545 8.515 3.55 ;
      RECT  7.3 3.55 8.515 3.555 ;
      RECT  7.305 3.555 8.515 3.56 ;
      RECT  7.31 3.56 8.515 3.565 ;
      RECT  7.315 3.565 8.515 3.57 ;
      RECT  7.32 3.57 8.515 3.575 ;
      RECT  7.325 3.575 8.515 3.58 ;
      RECT  7.33 3.58 8.515 3.585 ;
      RECT  7.335 3.585 8.515 3.59 ;
      RECT  7.34 3.59 8.515 3.595 ;
      RECT  7.345 3.595 8.515 3.6 ;
      RECT  7.35 3.6 8.515 3.605 ;
      RECT  7.355 3.605 8.515 3.61 ;
      RECT  7.36 3.61 8.515 3.615 ;
      RECT  7.365 3.615 8.515 3.62 ;
      RECT  7.37 3.62 8.515 3.625 ;
      RECT  7.375 3.625 8.515 3.63 ;
      RECT  7.38 3.63 8.515 3.635 ;
      RECT  7.385 3.635 8.515 3.64 ;
      RECT  7.39 3.64 8.515 3.645 ;
      RECT  7.395 3.645 8.515 3.65 ;
      RECT  7.4 3.65 8.515 3.655 ;
      RECT  7.405 3.655 8.515 3.66 ;
      RECT  7.41 3.66 8.515 3.665 ;
      RECT  7.415 3.665 8.515 3.67 ;
      RECT  7.42 3.67 8.515 3.675 ;
      RECT  7.425 3.675 8.515 3.68 ;
      RECT  7.43 3.68 8.515 3.685 ;
      RECT  7.435 3.685 8.515 3.69 ;
      RECT  7.44 3.69 8.515 3.695 ;
      RECT  7.445 3.695 8.515 3.7 ;
      RECT  7.45 3.7 8.515 3.705 ;
      RECT  7.455 3.705 8.515 3.71 ;
      RECT  7.46 3.71 8.515 3.715 ;
      RECT  7.465 3.715 8.515 3.72 ;
      RECT  7.47 3.72 8.515 3.725 ;
      RECT  7.475 3.725 8.515 3.73 ;
      RECT  7.48 3.73 8.515 3.735 ;
      RECT  7.485 3.735 8.515 3.74 ;
      RECT  7.49 3.74 8.515 3.745 ;
      RECT  7.495 3.745 8.515 3.75 ;
      RECT  7.5 3.75 8.515 3.755 ;
      RECT  7.505 3.755 8.515 3.76 ;
      RECT  7.51 3.76 8.515 3.765 ;
      RECT  7.515 3.765 8.515 3.77 ;
      RECT  7.52 3.77 8.515 3.775 ;
      RECT  2.42 3.62 5.0 3.85 ;
      RECT  2.125 4.08 4.3 4.31 ;
      RECT  2.125 4.31 2.355 4.365 ;
      RECT  0.18 4.365 2.355 4.595 ;
      RECT  5.025 4.62 6.175 4.85 ;
      RECT  5.025 4.85 5.255 5.0 ;
      RECT  5.945 4.85 6.175 5.0 ;
      RECT  3.75 5.0 5.255 5.23 ;
      RECT  5.945 5.0 7.45 5.23 ;
  END
END MDN_FDPQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPQ_2
#      Description : D-Flip Flop, pos-edge triggered, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPQ_2
  CLASS CORE ;
  FOREIGN MDN_FDPQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 4.365 11.9 5.0 ;
      RECT  11.59 5.0 11.93 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.92 1.565 13.96 1.795 ;
      RECT  13.325 1.795 13.555 3.245 ;
      RECT  12.92 3.245 13.96 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  5.485 5.08 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  5.48 1.005 6.22 1.235 ;
      RECT  5.48 1.235 5.71 1.565 ;
      RECT  3.19 1.565 5.71 1.795 ;
      RECT  4.36 1.795 4.59 3.03 ;
      RECT  3.19 3.03 4.59 3.26 ;
      RECT  10.47 0.37 10.81 0.6 ;
      RECT  10.47 0.6 10.7 1.005 ;
      RECT  7.725 1.005 10.7 1.235 ;
      RECT  7.725 1.235 7.955 3.315 ;
      RECT  12.71 0.37 14.17 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  10.975 1.005 12.94 1.235 ;
      RECT  10.975 1.235 11.205 1.565 ;
      RECT  10.525 1.565 11.205 1.795 ;
      RECT  10.525 1.795 10.755 2.405 ;
      RECT  9.35 2.405 10.755 2.635 ;
      RECT  10.525 2.635 10.755 3.245 ;
      RECT  10.525 3.245 11.02 3.475 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.005 5.0 1.235 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 2.38 ;
      RECT  2.685 2.38 4.09 2.61 ;
      RECT  2.685 2.61 2.915 3.03 ;
      RECT  1.72 3.03 2.915 3.26 ;
      RECT  6.045 1.565 7.24 1.795 ;
      RECT  6.045 1.795 6.275 2.405 ;
      RECT  4.87 2.405 6.275 2.635 ;
      RECT  6.045 2.635 6.275 3.7 ;
      RECT  6.045 3.7 7.095 3.93 ;
      RECT  6.865 3.93 7.095 4.005 ;
      RECT  6.865 4.005 8.78 4.235 ;
      RECT  8.44 1.565 9.48 1.795 ;
      RECT  11.435 1.51 11.875 1.85 ;
      RECT  11.645 1.85 11.875 3.805 ;
      RECT  9.405 3.805 11.875 4.035 ;
      RECT  9.405 4.035 9.635 5.0 ;
      RECT  4.53 4.16 6.635 4.39 ;
      RECT  4.53 4.39 4.76 4.465 ;
      RECT  6.405 4.39 6.635 4.465 ;
      RECT  2.74 4.465 4.76 4.695 ;
      RECT  6.405 4.465 8.46 4.695 ;
      RECT  2.74 4.695 2.97 5.0 ;
      RECT  8.23 4.695 8.46 5.0 ;
      RECT  1.51 5.0 2.97 5.23 ;
      RECT  8.23 5.0 9.635 5.23 ;
      RECT  8.285 3.245 9.48 3.475 ;
      RECT  8.285 3.475 8.515 3.545 ;
      RECT  6.9 3.24 7.325 3.245 ;
      RECT  6.9 3.245 7.33 3.25 ;
      RECT  6.9 3.25 7.335 3.255 ;
      RECT  6.9 3.255 7.34 3.26 ;
      RECT  6.9 3.26 7.345 3.265 ;
      RECT  6.9 3.265 7.35 3.27 ;
      RECT  6.9 3.27 7.355 3.275 ;
      RECT  6.9 3.275 7.36 3.28 ;
      RECT  6.9 3.28 7.365 3.285 ;
      RECT  6.9 3.285 7.37 3.29 ;
      RECT  6.9 3.29 7.375 3.295 ;
      RECT  6.9 3.295 7.38 3.3 ;
      RECT  6.9 3.3 7.385 3.305 ;
      RECT  6.9 3.305 7.39 3.31 ;
      RECT  6.9 3.31 7.395 3.315 ;
      RECT  6.9 3.315 7.4 3.32 ;
      RECT  6.9 3.32 7.405 3.325 ;
      RECT  6.9 3.325 7.41 3.33 ;
      RECT  6.9 3.33 7.415 3.335 ;
      RECT  6.9 3.335 7.42 3.34 ;
      RECT  6.9 3.34 7.425 3.345 ;
      RECT  6.9 3.345 7.43 3.35 ;
      RECT  6.9 3.35 7.435 3.355 ;
      RECT  6.9 3.355 7.44 3.36 ;
      RECT  6.9 3.36 7.445 3.365 ;
      RECT  6.9 3.365 7.45 3.37 ;
      RECT  6.9 3.37 7.455 3.375 ;
      RECT  6.9 3.375 7.46 3.38 ;
      RECT  6.9 3.38 7.465 3.385 ;
      RECT  6.9 3.385 7.47 3.39 ;
      RECT  6.9 3.39 7.475 3.395 ;
      RECT  6.9 3.395 7.48 3.4 ;
      RECT  6.9 3.4 7.485 3.405 ;
      RECT  6.9 3.405 7.49 3.41 ;
      RECT  6.9 3.41 7.495 3.415 ;
      RECT  6.9 3.415 7.5 3.42 ;
      RECT  6.9 3.42 7.505 3.425 ;
      RECT  6.9 3.425 7.51 3.43 ;
      RECT  6.9 3.43 7.515 3.435 ;
      RECT  6.9 3.435 7.52 3.44 ;
      RECT  6.9 3.44 7.525 3.445 ;
      RECT  6.9 3.445 7.53 3.45 ;
      RECT  6.9 3.45 7.535 3.455 ;
      RECT  6.9 3.455 7.54 3.46 ;
      RECT  6.9 3.46 7.545 3.465 ;
      RECT  6.9 3.465 7.55 3.47 ;
      RECT  7.22 3.47 7.555 3.475 ;
      RECT  7.225 3.475 7.56 3.48 ;
      RECT  7.23 3.48 7.565 3.485 ;
      RECT  7.235 3.485 7.57 3.49 ;
      RECT  7.24 3.49 7.575 3.495 ;
      RECT  7.245 3.495 7.58 3.5 ;
      RECT  7.25 3.5 7.585 3.505 ;
      RECT  7.255 3.505 7.59 3.51 ;
      RECT  7.26 3.51 7.595 3.515 ;
      RECT  7.265 3.515 7.6 3.52 ;
      RECT  7.27 3.52 7.605 3.525 ;
      RECT  7.275 3.525 7.61 3.53 ;
      RECT  7.28 3.53 7.615 3.535 ;
      RECT  7.285 3.535 7.62 3.54 ;
      RECT  7.29 3.54 7.625 3.545 ;
      RECT  7.295 3.545 8.515 3.55 ;
      RECT  7.3 3.55 8.515 3.555 ;
      RECT  7.305 3.555 8.515 3.56 ;
      RECT  7.31 3.56 8.515 3.565 ;
      RECT  7.315 3.565 8.515 3.57 ;
      RECT  7.32 3.57 8.515 3.575 ;
      RECT  7.325 3.575 8.515 3.58 ;
      RECT  7.33 3.58 8.515 3.585 ;
      RECT  7.335 3.585 8.515 3.59 ;
      RECT  7.34 3.59 8.515 3.595 ;
      RECT  7.345 3.595 8.515 3.6 ;
      RECT  7.35 3.6 8.515 3.605 ;
      RECT  7.355 3.605 8.515 3.61 ;
      RECT  7.36 3.61 8.515 3.615 ;
      RECT  7.365 3.615 8.515 3.62 ;
      RECT  7.37 3.62 8.515 3.625 ;
      RECT  7.375 3.625 8.515 3.63 ;
      RECT  7.38 3.63 8.515 3.635 ;
      RECT  7.385 3.635 8.515 3.64 ;
      RECT  7.39 3.64 8.515 3.645 ;
      RECT  7.395 3.645 8.515 3.65 ;
      RECT  7.4 3.65 8.515 3.655 ;
      RECT  7.405 3.655 8.515 3.66 ;
      RECT  7.41 3.66 8.515 3.665 ;
      RECT  7.415 3.665 8.515 3.67 ;
      RECT  7.42 3.67 8.515 3.675 ;
      RECT  7.425 3.675 8.515 3.68 ;
      RECT  7.43 3.68 8.515 3.685 ;
      RECT  7.435 3.685 8.515 3.69 ;
      RECT  7.44 3.69 8.515 3.695 ;
      RECT  7.445 3.695 8.515 3.7 ;
      RECT  7.45 3.7 8.515 3.705 ;
      RECT  7.455 3.705 8.515 3.71 ;
      RECT  7.46 3.71 8.515 3.715 ;
      RECT  7.465 3.715 8.515 3.72 ;
      RECT  7.47 3.72 8.515 3.725 ;
      RECT  7.475 3.725 8.515 3.73 ;
      RECT  7.48 3.73 8.515 3.735 ;
      RECT  7.485 3.735 8.515 3.74 ;
      RECT  7.49 3.74 8.515 3.745 ;
      RECT  7.495 3.745 8.515 3.75 ;
      RECT  7.5 3.75 8.515 3.755 ;
      RECT  7.505 3.755 8.515 3.76 ;
      RECT  7.51 3.76 8.515 3.765 ;
      RECT  7.515 3.765 8.515 3.77 ;
      RECT  7.52 3.77 8.515 3.775 ;
      RECT  2.42 3.51 5.0 3.74 ;
      RECT  2.125 3.98 4.3 4.21 ;
      RECT  2.125 4.21 2.355 4.365 ;
      RECT  0.18 4.365 2.355 4.595 ;
      RECT  5.025 4.62 6.175 4.85 ;
      RECT  5.025 4.85 5.255 4.925 ;
      RECT  5.945 4.85 6.175 5.0 ;
      RECT  3.75 4.925 5.255 5.155 ;
      RECT  5.945 5.0 7.45 5.23 ;
      RECT  3.75 5.155 4.09 5.23 ;
  END
END MDN_FDPQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPQ_4
#      Description : D-Flip Flop, pos-edge triggered, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPQ_4
  CLASS CORE ;
  FOREIGN MDN_FDPQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 4.365 11.9 5.0 ;
      RECT  11.59 5.0 11.93 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.92 1.565 16.2 1.795 ;
      RECT  14.445 1.795 14.675 3.245 ;
      RECT  12.92 3.245 16.2 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  5.485 5.08 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.66 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  5.485 1.005 6.22 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  3.19 1.565 5.715 1.795 ;
      RECT  4.365 1.795 4.595 3.16 ;
      RECT  3.19 3.16 4.595 3.39 ;
      RECT  10.425 0.37 10.81 0.6 ;
      RECT  10.425 0.6 10.655 1.005 ;
      RECT  7.745 1.005 10.655 1.235 ;
      RECT  7.745 1.235 7.975 3.315 ;
      RECT  14.95 0.37 16.41 0.6 ;
      RECT  14.95 0.6 15.18 1.005 ;
      RECT  12.71 0.37 14.17 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  13.94 0.6 14.17 1.005 ;
      RECT  10.885 1.005 12.94 1.235 ;
      RECT  13.94 1.005 15.18 1.235 ;
      RECT  10.885 1.235 11.115 1.565 ;
      RECT  10.525 1.565 11.115 1.795 ;
      RECT  10.525 1.795 10.755 2.405 ;
      RECT  9.35 2.405 10.755 2.635 ;
      RECT  10.525 2.635 10.755 3.17 ;
      RECT  10.525 3.17 11.02 3.4 ;
      RECT  0.14 1.005 2.76 1.235 ;
      RECT  3.96 1.005 5.0 1.235 ;
      RECT  1.72 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 2.395 ;
      RECT  2.125 2.395 3.95 2.625 ;
      RECT  2.125 2.625 2.355 3.165 ;
      RECT  1.72 3.165 2.355 3.395 ;
      RECT  6.045 1.565 7.24 1.795 ;
      RECT  6.045 1.795 6.275 2.405 ;
      RECT  4.87 2.405 6.275 2.635 ;
      RECT  6.045 2.635 6.275 3.7 ;
      RECT  6.045 3.7 7.095 3.93 ;
      RECT  6.865 3.93 7.095 4.015 ;
      RECT  6.865 4.015 8.78 4.245 ;
      RECT  8.44 1.565 9.48 1.795 ;
      RECT  11.38 1.565 11.875 1.795 ;
      RECT  11.645 1.795 11.875 3.805 ;
      RECT  9.405 3.805 11.875 4.035 ;
      RECT  9.405 4.035 9.635 4.475 ;
      RECT  4.565 4.16 6.635 4.39 ;
      RECT  6.405 4.39 6.635 4.475 ;
      RECT  4.565 4.39 4.795 4.54 ;
      RECT  6.405 4.475 9.635 4.705 ;
      RECT  2.76 4.54 4.795 4.77 ;
      RECT  8.23 4.705 8.46 5.0 ;
      RECT  2.76 4.77 2.99 5.0 ;
      RECT  1.51 5.0 2.99 5.23 ;
      RECT  8.23 5.0 8.57 5.23 ;
      RECT  8.285 3.245 9.48 3.475 ;
      RECT  8.285 3.475 8.515 3.545 ;
      RECT  6.9 3.24 7.345 3.245 ;
      RECT  6.9 3.245 7.35 3.25 ;
      RECT  6.9 3.25 7.355 3.255 ;
      RECT  6.9 3.255 7.36 3.26 ;
      RECT  6.9 3.26 7.365 3.265 ;
      RECT  6.9 3.265 7.37 3.27 ;
      RECT  6.9 3.27 7.375 3.275 ;
      RECT  6.9 3.275 7.38 3.28 ;
      RECT  6.9 3.28 7.385 3.285 ;
      RECT  6.9 3.285 7.39 3.29 ;
      RECT  6.9 3.29 7.395 3.295 ;
      RECT  6.9 3.295 7.4 3.3 ;
      RECT  6.9 3.3 7.405 3.305 ;
      RECT  6.9 3.305 7.41 3.31 ;
      RECT  6.9 3.31 7.415 3.315 ;
      RECT  6.9 3.315 7.42 3.32 ;
      RECT  6.9 3.32 7.425 3.325 ;
      RECT  6.9 3.325 7.43 3.33 ;
      RECT  6.9 3.33 7.435 3.335 ;
      RECT  6.9 3.335 7.44 3.34 ;
      RECT  6.9 3.34 7.445 3.345 ;
      RECT  6.9 3.345 7.45 3.35 ;
      RECT  6.9 3.35 7.455 3.355 ;
      RECT  6.9 3.355 7.46 3.36 ;
      RECT  6.9 3.36 7.465 3.365 ;
      RECT  6.9 3.365 7.47 3.37 ;
      RECT  6.9 3.37 7.475 3.375 ;
      RECT  6.9 3.375 7.48 3.38 ;
      RECT  6.9 3.38 7.485 3.385 ;
      RECT  6.9 3.385 7.49 3.39 ;
      RECT  6.9 3.39 7.495 3.395 ;
      RECT  6.9 3.395 7.5 3.4 ;
      RECT  6.9 3.4 7.505 3.405 ;
      RECT  6.9 3.405 7.51 3.41 ;
      RECT  6.9 3.41 7.515 3.415 ;
      RECT  6.9 3.415 7.52 3.42 ;
      RECT  6.9 3.42 7.525 3.425 ;
      RECT  6.9 3.425 7.53 3.43 ;
      RECT  6.9 3.43 7.535 3.435 ;
      RECT  6.9 3.435 7.54 3.44 ;
      RECT  6.9 3.44 7.545 3.445 ;
      RECT  6.9 3.445 7.55 3.45 ;
      RECT  6.9 3.45 7.555 3.455 ;
      RECT  6.9 3.455 7.56 3.46 ;
      RECT  6.9 3.46 7.565 3.465 ;
      RECT  6.9 3.465 7.57 3.47 ;
      RECT  7.24 3.47 7.575 3.475 ;
      RECT  7.245 3.475 7.58 3.48 ;
      RECT  7.25 3.48 7.585 3.485 ;
      RECT  7.255 3.485 7.59 3.49 ;
      RECT  7.26 3.49 7.595 3.495 ;
      RECT  7.265 3.495 7.6 3.5 ;
      RECT  7.27 3.5 7.605 3.505 ;
      RECT  7.275 3.505 7.61 3.51 ;
      RECT  7.28 3.51 7.615 3.515 ;
      RECT  7.285 3.515 7.62 3.52 ;
      RECT  7.29 3.52 7.625 3.525 ;
      RECT  7.295 3.525 7.63 3.53 ;
      RECT  7.3 3.53 7.635 3.535 ;
      RECT  7.305 3.535 7.64 3.54 ;
      RECT  7.31 3.54 7.645 3.545 ;
      RECT  7.315 3.545 8.515 3.55 ;
      RECT  7.32 3.55 8.515 3.555 ;
      RECT  7.325 3.555 8.515 3.56 ;
      RECT  7.33 3.56 8.515 3.565 ;
      RECT  7.335 3.565 8.515 3.57 ;
      RECT  7.34 3.57 8.515 3.575 ;
      RECT  7.345 3.575 8.515 3.58 ;
      RECT  7.35 3.58 8.515 3.585 ;
      RECT  7.355 3.585 8.515 3.59 ;
      RECT  7.36 3.59 8.515 3.595 ;
      RECT  7.365 3.595 8.515 3.6 ;
      RECT  7.37 3.6 8.515 3.605 ;
      RECT  7.375 3.605 8.515 3.61 ;
      RECT  7.38 3.61 8.515 3.615 ;
      RECT  7.385 3.615 8.515 3.62 ;
      RECT  7.39 3.62 8.515 3.625 ;
      RECT  7.395 3.625 8.515 3.63 ;
      RECT  7.4 3.63 8.515 3.635 ;
      RECT  7.405 3.635 8.515 3.64 ;
      RECT  7.41 3.64 8.515 3.645 ;
      RECT  7.415 3.645 8.515 3.65 ;
      RECT  7.42 3.65 8.515 3.655 ;
      RECT  7.425 3.655 8.515 3.66 ;
      RECT  7.43 3.66 8.515 3.665 ;
      RECT  7.435 3.665 8.515 3.67 ;
      RECT  7.44 3.67 8.515 3.675 ;
      RECT  7.445 3.675 8.515 3.68 ;
      RECT  7.45 3.68 8.515 3.685 ;
      RECT  7.455 3.685 8.515 3.69 ;
      RECT  7.46 3.69 8.515 3.695 ;
      RECT  7.465 3.695 8.515 3.7 ;
      RECT  7.47 3.7 8.515 3.705 ;
      RECT  7.475 3.705 8.515 3.71 ;
      RECT  7.48 3.71 8.515 3.715 ;
      RECT  7.485 3.715 8.515 3.72 ;
      RECT  7.49 3.72 8.515 3.725 ;
      RECT  7.495 3.725 8.515 3.73 ;
      RECT  7.5 3.73 8.515 3.735 ;
      RECT  7.505 3.735 8.515 3.74 ;
      RECT  7.51 3.74 8.515 3.745 ;
      RECT  7.515 3.745 8.515 3.75 ;
      RECT  7.52 3.75 8.515 3.755 ;
      RECT  7.525 3.755 8.515 3.76 ;
      RECT  7.53 3.76 8.515 3.765 ;
      RECT  7.535 3.765 8.515 3.77 ;
      RECT  7.54 3.77 8.515 3.775 ;
      RECT  2.42 3.62 5.0 3.85 ;
      RECT  2.125 4.08 4.3 4.31 ;
      RECT  2.125 4.31 2.355 4.365 ;
      RECT  0.14 4.365 2.355 4.595 ;
      RECT  5.025 4.62 6.175 4.85 ;
      RECT  5.025 4.85 5.255 5.0 ;
      RECT  5.945 4.85 6.175 5.0 ;
      RECT  3.75 5.0 5.255 5.23 ;
      RECT  5.945 5.0 7.45 5.23 ;
  END
END MDN_FDPQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPRB_4
#      Description : D-Flip Flop, pos-edge triggered, lo-async-clear
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPRB_4
  CLASS CORE ;
  FOREIGN MDN_FDPRB_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 24.64 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.16 1.565 18.44 1.795 ;
      RECT  17.805 1.795 18.035 3.245 ;
      RECT  15.16 3.245 18.445 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  20.33 1.565 24.46 1.795 ;
      RECT  22.285 1.795 22.515 3.245 ;
      RECT  20.34 3.245 24.46 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END QN
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 9.66 2.355 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.81 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  20.72 5.46 21.395 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  7.725 5.08 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 5.08 10.195 5.46 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 24.64 5.74 ;
      LAYER VIA12 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  24.23 5.47 24.49 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 -0.14 24.81 0.14 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  21.165 -0.14 21.84 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  16.685 -0.14 19.155 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  8.4 -0.14 9.52 0.14 ;
      RECT  8.845 0.14 9.075 0.89 ;
      RECT  8.44 0.89 9.48 1.12 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.6 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 24.64 0.14 ;
      LAYER VIA12 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  18.07 -0.13 18.33 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  9.965 0.37 11.93 0.6 ;
      RECT  9.965 0.6 10.195 1.35 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 0.83 ;
      RECT  1.565 0.83 6.22 1.005 ;
      RECT  1.565 1.005 7.955 1.06 ;
      RECT  1.565 1.06 2.06 1.12 ;
      RECT  5.99 1.06 7.955 1.235 ;
      RECT  1.565 1.12 1.795 3.805 ;
      RECT  7.725 1.235 7.955 1.35 ;
      RECT  7.725 1.35 10.195 1.58 ;
      RECT  1.565 3.805 2.06 4.035 ;
      RECT  19.43 0.37 19.77 0.6 ;
      RECT  19.43 0.6 19.66 1.005 ;
      RECT  17.19 0.37 18.65 0.6 ;
      RECT  18.42 0.6 18.65 1.005 ;
      RECT  18.42 1.005 19.66 1.235 ;
      RECT  21.67 0.37 23.13 0.6 ;
      RECT  10.68 1.005 14.675 1.235 ;
      RECT  14.445 1.235 14.675 2.125 ;
      RECT  13.885 2.125 17.475 2.355 ;
      RECT  15.005 2.355 15.235 2.69 ;
      RECT  16.125 2.355 16.355 2.69 ;
      RECT  17.245 2.355 17.475 2.69 ;
      RECT  13.885 2.355 14.115 4.02 ;
      RECT  9.14 4.02 14.115 4.25 ;
      RECT  2.42 1.29 5.0 1.52 ;
      RECT  5.43 1.565 5.77 1.795 ;
      RECT  5.43 1.795 5.66 2.405 ;
      RECT  3.75 2.405 5.66 2.635 ;
      RECT  5.43 2.635 5.66 3.03 ;
      RECT  5.43 3.03 5.77 3.26 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  10.525 1.565 11.72 1.795 ;
      RECT  10.525 1.795 10.755 1.81 ;
      RECT  9.965 1.81 10.755 2.04 ;
      RECT  9.965 2.04 10.195 3.49 ;
      RECT  3.245 1.75 4.3 1.98 ;
      RECT  3.245 1.98 3.475 3.49 ;
      RECT  3.245 3.49 13.26 3.72 ;
      RECT  7.165 2.35 7.395 3.49 ;
      RECT  12.15 1.565 12.49 1.795 ;
      RECT  12.15 1.795 12.38 2.405 ;
      RECT  10.47 2.405 12.38 2.635 ;
      RECT  12.15 2.635 12.38 3.03 ;
      RECT  12.15 3.03 12.49 3.26 ;
      RECT  12.92 1.565 13.96 1.795 ;
      RECT  19.485 1.565 19.98 1.795 ;
      RECT  19.485 1.795 19.715 2.125 ;
      RECT  19.485 2.125 21.955 2.355 ;
      RECT  20.605 2.355 20.835 2.69 ;
      RECT  21.725 2.355 21.955 2.69 ;
      RECT  19.485 2.355 19.715 3.245 ;
      RECT  19.485 3.245 19.98 3.475 ;
      RECT  22.845 2.125 24.195 2.355 ;
      RECT  22.845 2.355 23.075 2.69 ;
      RECT  23.965 2.355 24.195 2.69 ;
      RECT  2.42 3.95 6.54 4.18 ;
      RECT  6.805 4.1 8.78 4.33 ;
      RECT  6.805 4.33 7.035 4.41 ;
      RECT  4.66 4.41 7.035 4.64 ;
      RECT  11.38 4.48 13.96 4.71 ;
      RECT  7.265 4.56 10.755 4.79 ;
      RECT  7.265 4.79 7.495 5.0 ;
      RECT  10.525 4.79 10.755 5.0 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 1.74 4.41 ;
      RECT  0.18 4.41 4.035 4.595 ;
      RECT  1.51 4.595 4.035 4.64 ;
      RECT  1.51 4.64 1.74 5.0 ;
      RECT  3.805 4.64 4.035 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  3.805 5.0 7.495 5.23 ;
      RECT  10.525 5.0 13.05 5.23 ;
  END
END MDN_FDPRB_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPRB_1
#      Description : D-Flip Flop, pos-edge triggered, lo-async-clear
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPRB_1
  CLASS CORE ;
  FOREIGN MDN_FDPRB_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.86 1.565 16.915 1.795 ;
      RECT  16.685 1.795 16.915 3.245 ;
      RECT  15.86 3.245 16.915 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.245 1.565 17.74 1.795 ;
      RECT  17.245 1.795 17.475 3.245 ;
      RECT  17.245 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END QN
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.95 3.22 12.33 3.245 ;
      RECT  11.95 3.245 14.115 3.475 ;
      RECT  13.885 2.355 14.115 3.245 ;
      RECT  11.95 3.475 12.33 3.5 ;
      RECT  7.11 2.4 7.955 2.63 ;
      RECT  7.11 2.63 7.45 2.635 ;
      RECT  7.725 2.63 7.955 3.22 ;
      RECT  7.65 3.22 8.03 3.5 ;
      RECT  2.66 2.125 2.94 3.22 ;
      RECT  2.66 3.22 3.04 3.5 ;
      LAYER METAL2 ;
      RECT  2.66 3.22 12.33 3.5 ;
      LAYER VIA12 ;
      RECT  12.01 3.23 12.27 3.49 ;
      RECT  7.71 3.23 7.97 3.49 ;
      RECT  2.72 3.23 2.98 3.49 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  7.67 5.135 8.01 5.46 ;
      RECT  7.28 5.46 8.4 5.74 ;
      RECT  3.19 5.135 3.53 5.46 ;
      RECT  2.8 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  12.205 -0.14 14.115 0.14 ;
      RECT  12.205 0.14 12.435 0.6 ;
      RECT  13.885 0.14 14.115 0.89 ;
      RECT  13.62 0.89 14.115 1.12 ;
      RECT  6.72 -0.14 7.395 0.14 ;
      RECT  7.165 0.14 7.395 0.89 ;
      RECT  6.9 0.89 7.395 1.12 ;
      RECT  2.24 -0.14 2.915 0.14 ;
      RECT  2.685 0.14 2.915 1.005 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  9.02 0.37 11.93 0.38 ;
      RECT  9.01 0.38 11.93 0.6 ;
      RECT  9.01 0.6 9.24 1.225 ;
      RECT  9.005 1.225 9.24 1.23 ;
      RECT  9.0 1.23 9.24 1.235 ;
      RECT  8.995 1.235 9.24 1.24 ;
      RECT  8.99 1.24 9.24 1.245 ;
      RECT  8.985 1.245 9.24 1.25 ;
      RECT  8.98 1.25 9.24 1.255 ;
      RECT  8.975 1.255 9.24 1.26 ;
      RECT  8.97 1.26 9.24 1.265 ;
      RECT  8.965 1.265 9.24 1.27 ;
      RECT  8.96 1.27 9.24 1.275 ;
      RECT  8.955 1.275 9.24 1.28 ;
      RECT  8.95 1.28 9.24 1.285 ;
      RECT  8.945 1.285 9.24 1.29 ;
      RECT  8.94 1.29 9.24 1.295 ;
      RECT  8.935 1.295 9.24 1.3 ;
      RECT  8.93 1.3 9.24 1.305 ;
      RECT  8.925 1.305 9.24 1.31 ;
      RECT  8.92 1.31 9.24 1.315 ;
      RECT  8.915 1.315 9.24 1.32 ;
      RECT  8.91 1.32 9.235 1.325 ;
      RECT  8.905 1.325 9.23 1.33 ;
      RECT  8.9 1.33 9.225 1.335 ;
      RECT  8.895 1.335 9.22 1.34 ;
      RECT  8.89 1.34 9.215 1.345 ;
      RECT  8.885 1.345 9.21 1.35 ;
      RECT  8.88 1.35 9.205 1.355 ;
      RECT  8.875 1.355 9.2 1.36 ;
      RECT  8.87 1.36 9.195 1.365 ;
      RECT  8.865 1.365 9.19 1.37 ;
      RECT  8.86 1.37 9.185 1.375 ;
      RECT  8.855 1.375 9.18 1.38 ;
      RECT  8.85 1.38 9.175 1.385 ;
      RECT  8.845 1.385 9.17 1.39 ;
      RECT  8.84 1.39 9.165 1.395 ;
      RECT  8.835 1.395 9.16 1.4 ;
      RECT  8.83 1.4 9.155 1.405 ;
      RECT  8.825 1.405 9.15 1.41 ;
      RECT  8.82 1.41 9.145 1.415 ;
      RECT  8.815 1.415 9.14 1.42 ;
      RECT  8.81 1.42 9.135 1.425 ;
      RECT  8.805 1.425 9.13 1.43 ;
      RECT  8.8 1.43 9.125 1.435 ;
      RECT  8.795 1.435 9.12 1.44 ;
      RECT  8.79 1.44 9.115 1.445 ;
      RECT  8.785 1.445 9.11 1.45 ;
      RECT  8.78 1.45 9.105 1.455 ;
      RECT  8.775 1.455 9.1 1.46 ;
      RECT  8.77 1.46 9.095 1.465 ;
      RECT  8.765 1.465 9.09 1.47 ;
      RECT  8.76 1.47 9.085 1.475 ;
      RECT  8.755 1.475 9.08 1.48 ;
      RECT  8.75 1.48 9.075 1.485 ;
      RECT  8.745 1.485 9.07 1.49 ;
      RECT  8.74 1.49 9.065 1.495 ;
      RECT  8.735 1.495 9.06 1.5 ;
      RECT  8.73 1.5 9.055 1.505 ;
      RECT  8.725 1.505 9.05 1.51 ;
      RECT  8.72 1.51 9.045 1.515 ;
      RECT  8.715 1.515 9.04 1.52 ;
      RECT  8.71 1.52 9.035 1.525 ;
      RECT  8.705 1.525 9.03 1.53 ;
      RECT  8.7 1.53 9.025 1.535 ;
      RECT  8.695 1.535 9.02 1.54 ;
      RECT  8.69 1.54 9.015 1.545 ;
      RECT  8.685 1.545 9.01 1.55 ;
      RECT  8.68 1.55 9.005 1.555 ;
      RECT  8.675 1.555 9.0 1.56 ;
      RECT  8.67 1.56 8.995 1.565 ;
      RECT  8.665 1.565 8.99 1.57 ;
      RECT  8.66 1.57 8.985 1.575 ;
      RECT  8.655 1.575 8.98 1.58 ;
      RECT  8.65 1.58 8.975 1.585 ;
      RECT  8.645 1.585 8.97 1.59 ;
      RECT  8.64 1.59 8.965 1.595 ;
      RECT  8.635 1.595 8.96 1.6 ;
      RECT  8.63 1.6 8.955 1.605 ;
      RECT  8.625 1.605 8.95 1.61 ;
      RECT  8.62 1.61 8.945 1.615 ;
      RECT  8.615 1.615 8.94 1.62 ;
      RECT  8.61 1.62 8.935 1.625 ;
      RECT  8.605 1.625 8.93 1.63 ;
      RECT  8.6 1.63 8.925 1.635 ;
      RECT  8.595 1.635 8.92 1.64 ;
      RECT  8.59 1.64 8.915 1.645 ;
      RECT  8.585 1.645 8.91 1.65 ;
      RECT  8.58 1.65 8.905 1.655 ;
      RECT  8.575 1.655 8.9 1.66 ;
      RECT  8.57 1.66 8.895 1.665 ;
      RECT  8.565 1.665 8.89 1.67 ;
      RECT  8.56 1.67 8.885 1.675 ;
      RECT  8.555 1.675 8.88 1.68 ;
      RECT  8.55 1.68 8.875 1.685 ;
      RECT  8.545 1.685 8.87 1.69 ;
      RECT  8.54 1.69 8.865 1.695 ;
      RECT  8.535 1.695 8.86 1.7 ;
      RECT  8.53 1.7 8.855 1.705 ;
      RECT  8.525 1.705 8.85 1.71 ;
      RECT  8.52 1.71 8.845 1.715 ;
      RECT  8.515 1.715 8.84 1.72 ;
      RECT  8.51 1.72 8.835 1.725 ;
      RECT  8.505 1.725 8.83 1.73 ;
      RECT  8.5 1.73 8.825 1.735 ;
      RECT  8.495 1.735 8.82 1.74 ;
      RECT  8.49 1.74 8.815 1.745 ;
      RECT  8.485 1.745 8.81 1.75 ;
      RECT  8.48 1.75 8.805 1.755 ;
      RECT  8.475 1.755 8.8 1.76 ;
      RECT  8.47 1.76 8.795 1.765 ;
      RECT  8.465 1.765 8.79 1.77 ;
      RECT  8.46 1.77 8.785 1.775 ;
      RECT  8.455 1.775 8.78 1.78 ;
      RECT  8.45 1.78 8.775 1.785 ;
      RECT  8.445 1.785 8.77 1.79 ;
      RECT  8.44 1.79 8.765 1.795 ;
      RECT  8.435 1.795 8.76 1.8 ;
      RECT  8.43 1.8 8.755 1.805 ;
      RECT  8.425 1.805 8.75 1.81 ;
      RECT  5.38 1.75 5.72 1.81 ;
      RECT  5.38 1.81 8.745 1.815 ;
      RECT  5.38 1.815 8.74 1.82 ;
      RECT  5.38 1.82 8.735 1.825 ;
      RECT  5.38 1.825 8.73 1.83 ;
      RECT  5.38 1.83 8.725 1.835 ;
      RECT  5.38 1.835 8.72 1.84 ;
      RECT  5.38 1.84 8.715 1.845 ;
      RECT  5.38 1.845 8.71 1.85 ;
      RECT  5.38 1.85 8.705 1.855 ;
      RECT  5.38 1.855 8.7 1.86 ;
      RECT  5.38 1.86 8.695 1.865 ;
      RECT  5.38 1.865 8.69 1.87 ;
      RECT  5.38 1.87 8.685 1.875 ;
      RECT  5.38 1.875 8.68 1.88 ;
      RECT  5.38 1.88 8.675 1.885 ;
      RECT  5.38 1.885 8.67 1.89 ;
      RECT  5.38 1.89 8.665 1.895 ;
      RECT  5.38 1.895 8.66 1.9 ;
      RECT  5.38 1.9 8.655 1.905 ;
      RECT  5.38 1.905 8.65 1.91 ;
      RECT  5.38 1.91 8.645 1.915 ;
      RECT  5.38 1.915 8.64 1.92 ;
      RECT  5.38 1.92 8.635 1.925 ;
      RECT  5.38 1.925 8.63 1.93 ;
      RECT  5.38 1.93 8.625 1.935 ;
      RECT  5.38 1.935 8.62 1.94 ;
      RECT  5.38 1.94 8.615 1.945 ;
      RECT  5.38 1.945 8.61 1.95 ;
      RECT  5.38 1.95 8.605 1.955 ;
      RECT  5.38 1.955 8.6 1.96 ;
      RECT  5.38 1.96 8.595 1.965 ;
      RECT  5.38 1.965 8.59 1.97 ;
      RECT  5.38 1.97 8.585 1.975 ;
      RECT  5.38 1.975 8.58 1.98 ;
      RECT  5.38 1.98 8.575 1.985 ;
      RECT  5.38 1.985 8.57 1.99 ;
      RECT  5.38 1.99 8.565 1.995 ;
      RECT  5.38 1.995 8.56 2.0 ;
      RECT  5.38 2.0 8.555 2.005 ;
      RECT  5.38 2.005 8.55 2.01 ;
      RECT  5.38 2.01 8.545 2.015 ;
      RECT  5.38 2.015 8.54 2.02 ;
      RECT  5.38 2.02 8.535 2.025 ;
      RECT  5.38 2.025 8.53 2.03 ;
      RECT  5.38 2.03 8.525 2.035 ;
      RECT  5.38 2.035 8.52 2.04 ;
      RECT  6.605 2.04 6.835 3.245 ;
      RECT  5.43 3.245 7.24 3.475 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 1.74 1.235 ;
      RECT  3.245 0.37 5.21 0.6 ;
      RECT  3.245 0.6 3.475 1.565 ;
      RECT  1.005 1.565 3.475 1.795 ;
      RECT  1.005 1.795 1.235 3.805 ;
      RECT  1.005 3.805 2.355 4.035 ;
      RECT  2.125 4.035 2.355 4.215 ;
      RECT  2.125 4.215 10.195 4.445 ;
      RECT  9.965 4.445 10.195 5.0 ;
      RECT  9.965 5.0 10.81 5.23 ;
      RECT  17.19 0.37 17.53 0.6 ;
      RECT  17.19 0.6 17.42 1.005 ;
      RECT  14.445 0.37 16.355 0.6 ;
      RECT  16.125 0.6 16.355 1.005 ;
      RECT  14.445 0.6 14.675 1.35 ;
      RECT  16.125 1.005 17.42 1.235 ;
      RECT  9.965 1.29 12.45 1.35 ;
      RECT  9.965 1.35 14.675 1.52 ;
      RECT  12.18 1.52 14.675 1.58 ;
      RECT  9.965 1.52 10.195 3.465 ;
      RECT  4.015 0.83 6.54 1.06 ;
      RECT  6.2 1.06 6.54 1.12 ;
      RECT  4.015 1.06 4.245 1.29 ;
      RECT  9.475 0.83 13.26 1.06 ;
      RECT  12.92 1.06 13.26 1.12 ;
      RECT  9.475 1.06 9.705 1.75 ;
      RECT  9.14 1.75 9.705 1.98 ;
      RECT  7.725 0.89 8.78 1.12 ;
      RECT  7.725 1.12 7.955 1.35 ;
      RECT  4.66 1.29 6.045 1.35 ;
      RECT  4.66 1.35 7.955 1.52 ;
      RECT  5.875 1.52 7.955 1.58 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 1.895 ;
      RECT  12.765 1.895 15.235 2.125 ;
      RECT  12.765 2.125 12.995 2.62 ;
      RECT  15.005 2.125 15.235 2.685 ;
      RECT  15.005 2.685 16.355 2.915 ;
      RECT  16.125 2.35 16.355 2.685 ;
      RECT  15.005 2.915 15.235 3.805 ;
      RECT  13.62 3.805 15.5 4.035 ;
      RECT  10.68 1.75 11.72 1.98 ;
      RECT  11.085 1.98 11.315 3.245 ;
      RECT  11.085 3.245 11.72 3.475 ;
      RECT  11.085 3.475 11.315 3.705 ;
      RECT  8.23 2.405 9.36 2.635 ;
      RECT  9.13 2.635 9.36 3.705 ;
      RECT  9.13 3.705 11.315 3.935 ;
      RECT  3.96 3.245 5.0 3.475 ;
      RECT  6.2 3.755 8.78 3.985 ;
      RECT  0.18 4.365 1.85 4.595 ;
      RECT  1.62 4.595 1.85 4.675 ;
      RECT  1.62 4.675 9.58 4.905 ;
      RECT  1.62 4.905 1.85 5.0 ;
      RECT  9.35 4.905 9.58 5.0 ;
      RECT  5.99 4.905 6.33 5.23 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  9.35 5.0 9.69 5.23 ;
      RECT  10.68 4.365 13.26 4.595 ;
  END
END MDN_FDPRB_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPRB_2
#      Description : D-Flip Flop, pos-edge triggered, lo-async-clear
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPRB_2
  CLASS CORE ;
  FOREIGN MDN_FDPRB_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.86 1.565 17.74 1.795 ;
      RECT  16.685 1.795 16.915 3.245 ;
      RECT  15.86 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.1 1.565 19.98 1.795 ;
      RECT  18.925 1.795 19.155 3.245 ;
      RECT  18.1 3.245 19.98 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END QN
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.01 3.22 11.39 3.245 ;
      RECT  11.01 3.245 14.115 3.475 ;
      RECT  13.885 2.35 14.115 3.245 ;
      RECT  11.01 3.475 11.39 3.5 ;
      RECT  7.165 2.35 7.395 2.685 ;
      RECT  7.165 2.685 7.955 2.915 ;
      RECT  7.725 2.915 7.955 3.245 ;
      RECT  7.725 3.245 8.91 3.475 ;
      RECT  8.53 3.22 8.91 3.245 ;
      RECT  8.53 3.475 8.91 3.5 ;
      RECT  2.66 2.35 2.94 3.22 ;
      RECT  2.66 3.22 3.04 3.5 ;
      LAYER METAL2 ;
      RECT  2.66 3.22 11.39 3.5 ;
      LAYER VIA12 ;
      RECT  11.07 3.23 11.33 3.49 ;
      RECT  8.59 3.23 8.85 3.49 ;
      RECT  2.72 3.23 2.98 3.49 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  14.445 4.87 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  7.67 5.135 8.01 5.46 ;
      RECT  7.28 5.46 9.13 5.74 ;
      RECT  3.19 5.135 3.53 5.46 ;
      RECT  2.8 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  12.205 -0.14 14.115 0.14 ;
      RECT  12.205 0.14 12.435 0.6 ;
      RECT  13.885 0.14 14.115 0.89 ;
      RECT  13.62 0.89 14.115 1.12 ;
      RECT  6.72 -0.14 7.395 0.14 ;
      RECT  7.165 0.14 7.395 0.89 ;
      RECT  6.9 0.89 7.395 1.12 ;
      RECT  2.24 -0.14 2.915 0.14 ;
      RECT  2.685 0.14 2.915 1.005 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 1.74 1.235 ;
      RECT  3.245 0.37 5.21 0.6 ;
      RECT  3.245 0.6 3.475 1.565 ;
      RECT  1.005 1.565 3.475 1.795 ;
      RECT  1.005 1.795 1.235 3.805 ;
      RECT  1.005 3.805 2.355 4.035 ;
      RECT  2.125 4.035 2.355 4.215 ;
      RECT  2.125 4.215 10.195 4.445 ;
      RECT  9.965 4.445 10.195 5.0 ;
      RECT  9.965 5.0 10.81 5.23 ;
      RECT  9.01 0.37 11.93 0.6 ;
      RECT  9.01 0.6 9.24 1.225 ;
      RECT  9.005 1.225 9.24 1.23 ;
      RECT  9.0 1.23 9.24 1.235 ;
      RECT  8.995 1.235 9.24 1.24 ;
      RECT  8.99 1.24 9.24 1.245 ;
      RECT  8.985 1.245 9.24 1.25 ;
      RECT  8.98 1.25 9.24 1.255 ;
      RECT  8.975 1.255 9.24 1.26 ;
      RECT  8.97 1.26 9.24 1.265 ;
      RECT  8.965 1.265 9.24 1.27 ;
      RECT  8.96 1.27 9.24 1.275 ;
      RECT  8.955 1.275 9.24 1.28 ;
      RECT  8.95 1.28 9.24 1.285 ;
      RECT  8.945 1.285 9.24 1.29 ;
      RECT  8.94 1.29 9.24 1.295 ;
      RECT  8.935 1.295 9.24 1.3 ;
      RECT  8.93 1.3 9.24 1.305 ;
      RECT  8.925 1.305 9.24 1.31 ;
      RECT  8.92 1.31 9.24 1.315 ;
      RECT  8.915 1.315 9.24 1.32 ;
      RECT  8.91 1.32 9.235 1.325 ;
      RECT  8.905 1.325 9.23 1.33 ;
      RECT  8.9 1.33 9.225 1.335 ;
      RECT  8.895 1.335 9.22 1.34 ;
      RECT  8.89 1.34 9.215 1.345 ;
      RECT  8.885 1.345 9.21 1.35 ;
      RECT  8.285 1.35 9.205 1.355 ;
      RECT  8.285 1.355 9.2 1.36 ;
      RECT  8.285 1.36 9.195 1.365 ;
      RECT  8.285 1.365 9.19 1.37 ;
      RECT  8.285 1.37 9.185 1.375 ;
      RECT  8.285 1.375 9.18 1.38 ;
      RECT  8.285 1.38 9.175 1.385 ;
      RECT  8.285 1.385 9.17 1.39 ;
      RECT  8.285 1.39 9.165 1.395 ;
      RECT  8.285 1.395 9.16 1.4 ;
      RECT  8.285 1.4 9.155 1.405 ;
      RECT  8.285 1.405 9.15 1.41 ;
      RECT  8.285 1.41 9.145 1.415 ;
      RECT  8.285 1.415 9.14 1.42 ;
      RECT  8.285 1.42 9.135 1.425 ;
      RECT  8.285 1.425 9.13 1.43 ;
      RECT  8.285 1.43 9.125 1.435 ;
      RECT  8.285 1.435 9.12 1.44 ;
      RECT  8.285 1.44 9.115 1.445 ;
      RECT  8.285 1.445 9.11 1.45 ;
      RECT  8.285 1.45 9.105 1.455 ;
      RECT  8.285 1.455 9.1 1.46 ;
      RECT  8.285 1.46 9.095 1.465 ;
      RECT  8.285 1.465 9.09 1.47 ;
      RECT  8.285 1.47 9.085 1.475 ;
      RECT  8.285 1.475 9.08 1.48 ;
      RECT  8.285 1.48 9.075 1.485 ;
      RECT  8.285 1.485 9.07 1.49 ;
      RECT  8.285 1.49 9.065 1.495 ;
      RECT  8.285 1.495 9.06 1.5 ;
      RECT  8.285 1.5 9.055 1.505 ;
      RECT  8.285 1.505 9.05 1.51 ;
      RECT  8.285 1.51 9.045 1.515 ;
      RECT  8.285 1.515 9.04 1.52 ;
      RECT  8.285 1.52 9.035 1.525 ;
      RECT  8.285 1.525 9.03 1.53 ;
      RECT  8.285 1.53 9.025 1.535 ;
      RECT  8.285 1.535 9.02 1.54 ;
      RECT  8.285 1.54 9.015 1.545 ;
      RECT  8.285 1.545 9.01 1.55 ;
      RECT  8.285 1.55 9.005 1.555 ;
      RECT  8.285 1.555 9.0 1.56 ;
      RECT  8.285 1.56 8.995 1.565 ;
      RECT  8.285 1.565 8.99 1.57 ;
      RECT  8.285 1.57 8.985 1.575 ;
      RECT  8.285 1.575 8.98 1.58 ;
      RECT  8.285 1.58 8.515 1.81 ;
      RECT  5.43 1.75 5.77 1.81 ;
      RECT  5.43 1.81 8.515 2.04 ;
      RECT  6.605 2.04 6.835 3.17 ;
      RECT  5.43 3.17 7.24 3.4 ;
      RECT  19.43 0.37 19.77 0.6 ;
      RECT  19.43 0.6 19.66 1.005 ;
      RECT  18.31 0.37 18.65 0.6 ;
      RECT  18.42 0.6 18.65 1.005 ;
      RECT  14.445 0.37 16.355 0.6 ;
      RECT  16.125 0.6 16.355 1.005 ;
      RECT  14.445 0.6 14.675 1.35 ;
      RECT  16.125 1.005 19.66 1.235 ;
      RECT  9.965 1.29 12.435 1.35 ;
      RECT  9.965 1.35 14.675 1.52 ;
      RECT  12.205 1.52 14.675 1.58 ;
      RECT  9.965 1.52 10.195 3.46 ;
      RECT  3.96 0.83 6.54 1.06 ;
      RECT  6.2 1.06 6.54 1.12 ;
      RECT  3.96 1.06 4.3 1.235 ;
      RECT  9.47 0.83 13.26 1.06 ;
      RECT  12.92 1.06 13.26 1.12 ;
      RECT  9.47 1.06 9.7 1.75 ;
      RECT  9.14 1.75 9.7 1.98 ;
      RECT  7.725 0.89 8.78 1.12 ;
      RECT  7.725 1.12 7.955 1.35 ;
      RECT  4.715 1.29 5.98 1.295 ;
      RECT  4.715 1.295 5.985 1.3 ;
      RECT  4.715 1.3 5.99 1.305 ;
      RECT  4.715 1.305 5.995 1.31 ;
      RECT  4.715 1.31 6.0 1.315 ;
      RECT  4.715 1.315 6.005 1.32 ;
      RECT  4.715 1.32 6.01 1.325 ;
      RECT  4.715 1.325 6.015 1.33 ;
      RECT  4.715 1.33 6.02 1.335 ;
      RECT  4.715 1.335 6.025 1.34 ;
      RECT  4.715 1.34 6.03 1.345 ;
      RECT  4.715 1.345 6.035 1.35 ;
      RECT  4.715 1.35 7.955 1.52 ;
      RECT  5.875 1.52 7.955 1.525 ;
      RECT  4.715 1.52 4.945 1.85 ;
      RECT  5.88 1.525 7.955 1.53 ;
      RECT  5.885 1.53 7.955 1.535 ;
      RECT  5.89 1.535 7.955 1.54 ;
      RECT  5.895 1.54 7.955 1.545 ;
      RECT  5.9 1.545 7.955 1.55 ;
      RECT  5.905 1.55 7.955 1.555 ;
      RECT  5.91 1.555 7.955 1.56 ;
      RECT  5.915 1.56 7.955 1.565 ;
      RECT  5.92 1.565 7.955 1.57 ;
      RECT  5.925 1.57 7.955 1.575 ;
      RECT  5.93 1.575 7.955 1.58 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 1.81 ;
      RECT  12.765 1.81 15.235 2.04 ;
      RECT  12.765 2.04 12.995 2.69 ;
      RECT  15.005 2.04 15.235 4.365 ;
      RECT  13.62 4.365 17.42 4.595 ;
      RECT  16.18 4.595 16.41 5.0 ;
      RECT  17.19 4.595 17.42 5.0 ;
      RECT  16.07 5.0 16.41 5.23 ;
      RECT  17.19 5.0 17.53 5.23 ;
      RECT  10.525 1.75 11.72 1.98 ;
      RECT  10.525 1.98 10.755 3.755 ;
      RECT  8.23 2.405 9.635 2.635 ;
      RECT  9.405 2.635 9.635 3.245 ;
      RECT  9.14 3.245 9.635 3.475 ;
      RECT  9.405 3.475 9.635 3.755 ;
      RECT  9.405 3.755 11.72 3.985 ;
      RECT  3.96 3.755 5.0 3.985 ;
      RECT  6.2 3.755 8.78 3.985 ;
      RECT  0.18 4.365 1.85 4.595 ;
      RECT  1.51 4.595 1.85 4.675 ;
      RECT  1.51 4.675 9.475 4.905 ;
      RECT  9.245 4.905 9.475 5.0 ;
      RECT  1.51 4.905 1.85 5.23 ;
      RECT  5.99 4.905 6.33 5.23 ;
      RECT  9.245 5.0 9.69 5.23 ;
      RECT  10.68 4.365 13.26 4.595 ;
  END
END MDN_FDPRB_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPRBQ_F_1
#      Description : D-Flip Flop, pos-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPRBQ_F_1
  CLASS CORE ;
  FOREIGN MDN_FDPRBQ_F_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.98 0.37 1.85 0.6 ;
      RECT  0.98 0.6 1.26 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.245 1.565 17.74 1.795 ;
      RECT  17.245 1.795 17.475 3.245 ;
      RECT  17.245 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.97 4.545 15.16 4.775 ;
      RECT  13.97 4.775 14.2 4.925 ;
      RECT  14.93 4.775 15.16 5.0 ;
      RECT  7.725 4.365 10.755 4.535 ;
      RECT  7.24 4.535 10.755 4.595 ;
      RECT  7.24 4.595 8.44 4.765 ;
      RECT  10.525 4.595 10.755 4.925 ;
      RECT  7.24 4.765 7.47 4.925 ;
      RECT  8.21 4.765 8.44 5.0 ;
      RECT  0.42 4.365 3.965 4.595 ;
      RECT  3.55 4.595 3.965 4.62 ;
      RECT  0.42 4.595 0.7 5.0 ;
      RECT  3.735 4.62 3.965 4.925 ;
      RECT  3.735 4.925 7.47 5.155 ;
      RECT  10.525 4.925 14.2 5.155 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  8.21 5.0 8.57 5.23 ;
      RECT  14.93 5.0 15.29 5.23 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 5.005 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  7.725 4.995 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 4.995 10.195 5.46 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.56 -0.14 15.235 0.14 ;
      RECT  15.005 0.14 15.235 1.005 ;
      RECT  15.005 1.005 15.5 1.235 ;
      RECT  8.285 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.57 ;
      RECT  8.285 0.14 8.515 1.005 ;
      RECT  8.285 1.005 8.78 1.235 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 10.81 0.6 ;
      RECT  10.47 0.6 10.7 0.8 ;
      RECT  9.195 0.8 10.7 1.03 ;
      RECT  9.195 1.03 9.425 1.29 ;
      RECT  11.085 0.37 13.05 0.6 ;
      RECT  11.085 0.6 11.315 1.26 ;
      RECT  9.965 1.26 11.315 1.49 ;
      RECT  9.965 1.49 10.195 1.52 ;
      RECT  3.75 0.37 7.955 0.6 ;
      RECT  7.725 0.6 7.955 1.52 ;
      RECT  7.725 1.52 10.195 1.75 ;
      RECT  1.72 1.005 5.0 1.235 ;
      RECT  6.2 1.005 7.24 1.235 ;
      RECT  12.92 1.005 13.96 1.235 ;
      RECT  12.15 1.465 13.555 1.695 ;
      RECT  13.325 1.695 13.555 2.71 ;
      RECT  13.325 2.71 13.72 2.94 ;
      RECT  13.49 2.94 13.72 3.625 ;
      RECT  12.205 3.625 16.41 3.855 ;
      RECT  12.205 3.855 12.435 4.09 ;
      RECT  16.18 3.855 16.41 4.365 ;
      RECT  16.18 4.365 17.42 4.595 ;
      RECT  16.18 4.595 16.41 5.0 ;
      RECT  17.19 4.595 17.42 5.0 ;
      RECT  16.07 5.0 16.41 5.23 ;
      RECT  17.19 5.0 17.53 5.23 ;
      RECT  2.42 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 2.405 ;
      RECT  3.245 2.405 4.09 2.635 ;
      RECT  3.245 2.635 3.475 3.245 ;
      RECT  2.42 3.245 3.475 3.475 ;
      RECT  3.955 1.565 5.095 1.795 ;
      RECT  4.865 1.795 5.095 3.03 ;
      RECT  3.96 3.03 5.095 3.26 ;
      RECT  4.865 3.26 5.095 3.545 ;
      RECT  4.865 3.545 11.875 3.775 ;
      RECT  6.045 2.35 6.275 3.545 ;
      RECT  11.645 2.39 11.875 3.545 ;
      RECT  14.075 1.565 16.2 1.795 ;
      RECT  14.075 1.795 14.305 3.1 ;
      RECT  14.075 3.1 16.2 3.33 ;
      RECT  10.68 1.72 11.72 1.93 ;
      RECT  10.68 1.93 12.435 1.95 ;
      RECT  11.085 1.95 12.435 2.16 ;
      RECT  11.085 2.16 11.315 3.03 ;
      RECT  12.205 2.16 12.435 3.165 ;
      RECT  10.68 3.03 11.315 3.26 ;
      RECT  12.205 3.165 13.26 3.395 ;
      RECT  7.165 1.98 10.195 2.21 ;
      RECT  9.965 2.21 10.195 2.41 ;
      RECT  7.165 2.21 7.395 2.71 ;
      RECT  9.965 2.41 10.81 2.64 ;
      RECT  9.965 2.64 10.195 3.03 ;
      RECT  9.14 3.03 10.195 3.26 ;
      RECT  8.55 2.445 9.69 2.675 ;
      RECT  8.55 2.675 8.78 3.03 ;
      RECT  5.485 1.565 6.835 1.795 ;
      RECT  6.605 1.795 6.835 3.03 ;
      RECT  5.485 1.795 5.715 3.315 ;
      RECT  6.605 3.03 8.78 3.26 ;
      RECT  1.72 3.805 4.425 4.035 ;
      RECT  4.195 4.035 4.425 4.465 ;
      RECT  4.195 4.465 6.54 4.695 ;
      RECT  4.66 4.005 7.24 4.235 ;
      RECT  13.325 4.085 15.5 4.315 ;
      RECT  13.325 4.315 13.555 4.365 ;
      RECT  11.38 4.365 13.555 4.595 ;
  END
END MDN_FDPRBQ_F_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPRBQ_F_2
#      Description : D-Flip Flop, pos-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPRBQ_F_2
  CLASS CORE ;
  FOREIGN MDN_FDPRBQ_F_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.98 0.37 1.85 0.6 ;
      RECT  0.98 0.6 1.26 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.4 1.565 19.155 1.795 ;
      RECT  18.925 1.795 19.155 3.245 ;
      RECT  17.4 3.245 19.155 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.97 4.55 15.16 4.78 ;
      RECT  13.97 4.78 14.2 4.925 ;
      RECT  14.93 4.78 15.16 5.0 ;
      RECT  7.15 4.41 10.755 4.64 ;
      RECT  7.15 4.64 7.38 4.925 ;
      RECT  10.525 4.64 10.755 4.925 ;
      RECT  8.22 4.64 8.45 5.0 ;
      RECT  0.42 4.365 3.97 4.595 ;
      RECT  3.55 4.595 3.97 4.62 ;
      RECT  0.42 4.595 0.7 5.0 ;
      RECT  3.74 4.62 3.97 4.925 ;
      RECT  3.74 4.925 7.38 5.155 ;
      RECT  10.525 4.925 14.2 5.155 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  8.22 5.0 8.57 5.23 ;
      RECT  14.93 5.0 15.29 5.23 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  14.445 5.01 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.56 -0.14 15.235 0.14 ;
      RECT  15.005 0.14 15.235 1.005 ;
      RECT  15.005 1.005 15.5 1.235 ;
      RECT  8.285 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.57 ;
      RECT  8.285 0.14 8.515 1.005 ;
      RECT  8.285 1.005 8.78 1.235 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  12.71 0.37 13.05 0.445 ;
      RECT  11.085 0.445 13.05 0.675 ;
      RECT  11.085 0.675 11.315 1.26 ;
      RECT  9.94 1.26 11.315 1.465 ;
      RECT  3.75 0.37 7.955 0.6 ;
      RECT  7.725 0.6 7.955 1.465 ;
      RECT  7.725 1.465 11.315 1.49 ;
      RECT  7.725 1.49 10.17 1.695 ;
      RECT  10.47 0.37 10.81 0.6 ;
      RECT  10.47 0.6 10.7 0.8 ;
      RECT  9.14 0.8 10.7 1.03 ;
      RECT  9.14 1.03 9.48 1.235 ;
      RECT  1.72 1.005 5.0 1.235 ;
      RECT  6.2 1.005 7.24 1.235 ;
      RECT  12.92 1.005 13.96 1.235 ;
      RECT  2.42 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 2.405 ;
      RECT  3.245 2.405 4.09 2.635 ;
      RECT  3.245 2.635 3.475 3.245 ;
      RECT  2.42 3.245 3.475 3.475 ;
      RECT  14.075 1.565 16.2 1.795 ;
      RECT  14.075 1.795 14.305 3.03 ;
      RECT  14.075 3.03 16.2 3.26 ;
      RECT  10.68 1.72 11.72 1.935 ;
      RECT  10.68 1.935 12.435 1.95 ;
      RECT  11.085 1.95 12.435 2.165 ;
      RECT  11.085 2.165 11.315 3.03 ;
      RECT  12.205 2.165 12.435 3.03 ;
      RECT  10.735 3.03 11.315 3.26 ;
      RECT  12.205 3.03 13.26 3.26 ;
      RECT  10.735 3.26 10.965 3.53 ;
      RECT  7.165 1.925 10.195 2.155 ;
      RECT  9.965 2.155 10.195 2.445 ;
      RECT  7.165 2.155 7.395 2.69 ;
      RECT  9.965 2.445 10.81 2.675 ;
      RECT  9.965 2.675 10.195 3.03 ;
      RECT  9.195 3.03 10.195 3.26 ;
      RECT  9.195 3.26 9.425 3.53 ;
      RECT  9.35 2.445 9.69 2.475 ;
      RECT  8.495 2.475 9.69 2.705 ;
      RECT  8.495 2.705 8.725 3.03 ;
      RECT  5.485 1.695 6.835 1.925 ;
      RECT  5.485 1.925 5.715 3.03 ;
      RECT  6.605 1.925 6.835 3.03 ;
      RECT  5.43 3.03 5.77 3.26 ;
      RECT  6.605 3.03 8.725 3.26 ;
      RECT  8.495 3.26 8.725 3.53 ;
      RECT  11.59 2.405 11.93 2.635 ;
      RECT  11.645 2.635 11.875 3.805 ;
      RECT  3.955 1.565 4.595 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  3.96 3.245 5.155 3.475 ;
      RECT  4.925 3.475 5.155 3.49 ;
      RECT  4.925 3.49 7.985 3.72 ;
      RECT  6.045 2.35 6.275 3.49 ;
      RECT  7.755 3.72 7.985 3.805 ;
      RECT  7.755 3.805 11.875 4.035 ;
      RECT  16.07 2.405 18.43 2.635 ;
      RECT  16.685 2.635 16.915 3.49 ;
      RECT  12.15 1.475 13.72 1.705 ;
      RECT  13.49 1.705 13.72 3.49 ;
      RECT  12.205 3.49 16.915 3.72 ;
      RECT  12.205 3.72 12.435 4.09 ;
      RECT  1.72 3.805 4.43 4.035 ;
      RECT  4.2 4.035 4.43 4.41 ;
      RECT  4.2 4.41 6.54 4.64 ;
      RECT  4.66 3.95 7.24 4.18 ;
      RECT  13.325 4.09 15.5 4.32 ;
      RECT  13.325 4.32 13.555 4.365 ;
      RECT  11.38 4.365 13.555 4.595 ;
  END
END MDN_FDPRBQ_F_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPRBQ_F_4
#      Description : D-Flip Flop, pos-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPRBQ_F_4
  CLASS CORE ;
  FOREIGN MDN_FDPRBQ_F_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.98 0.37 1.85 0.6 ;
      RECT  0.98 0.6 1.26 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.4 1.565 21.395 1.795 ;
      RECT  21.165 1.795 21.395 3.245 ;
      RECT  17.4 3.245 21.395 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.96 4.55 15.16 4.78 ;
      RECT  13.96 4.78 14.19 4.925 ;
      RECT  14.93 4.78 15.16 5.0 ;
      RECT  7.725 4.365 10.755 4.465 ;
      RECT  7.24 4.465 10.755 4.595 ;
      RECT  7.24 4.595 8.44 4.695 ;
      RECT  10.525 4.595 10.755 4.925 ;
      RECT  7.24 4.695 7.47 4.925 ;
      RECT  8.21 4.695 8.44 5.0 ;
      RECT  0.42 4.365 3.935 4.595 ;
      RECT  3.55 4.595 3.935 4.62 ;
      RECT  0.42 4.595 0.7 5.0 ;
      RECT  3.705 4.62 3.935 4.925 ;
      RECT  3.705 4.925 7.47 5.155 ;
      RECT  10.525 4.925 14.19 5.155 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  8.21 5.0 8.57 5.23 ;
      RECT  14.93 5.0 15.29 5.23 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.925 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.925 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.925 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  14.445 5.01 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  7.725 4.93 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.925 -0.14 19.6 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.56 -0.14 15.235 0.14 ;
      RECT  15.005 0.14 15.235 1.005 ;
      RECT  15.005 1.005 15.5 1.235 ;
      RECT  8.285 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.57 ;
      RECT  8.285 0.14 8.515 1.005 ;
      RECT  8.285 1.005 8.78 1.235 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  12.71 0.37 13.05 0.445 ;
      RECT  11.085 0.445 13.05 0.675 ;
      RECT  11.085 0.675 11.315 1.26 ;
      RECT  9.965 1.26 11.315 1.49 ;
      RECT  9.965 1.49 10.195 1.52 ;
      RECT  3.75 0.37 7.955 0.6 ;
      RECT  7.725 0.6 7.955 1.52 ;
      RECT  7.725 1.52 10.195 1.75 ;
      RECT  10.47 0.37 10.81 0.6 ;
      RECT  10.47 0.6 10.7 0.8 ;
      RECT  9.195 0.8 10.7 1.03 ;
      RECT  9.195 1.03 9.425 1.29 ;
      RECT  1.72 1.005 5.0 1.235 ;
      RECT  6.2 1.005 7.24 1.235 ;
      RECT  12.92 1.005 13.96 1.235 ;
      RECT  2.42 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 2.415 ;
      RECT  3.245 2.415 4.09 2.645 ;
      RECT  3.245 2.645 3.475 3.245 ;
      RECT  2.42 3.245 3.475 3.475 ;
      RECT  3.955 1.565 4.595 1.795 ;
      RECT  4.365 1.795 4.595 3.03 ;
      RECT  3.96 3.03 5.155 3.26 ;
      RECT  4.925 3.26 5.155 3.545 ;
      RECT  4.925 3.545 11.875 3.775 ;
      RECT  6.045 2.35 6.275 3.545 ;
      RECT  11.645 2.39 11.875 3.545 ;
      RECT  15.565 1.565 16.2 1.795 ;
      RECT  15.565 1.795 15.795 2.335 ;
      RECT  14.01 2.335 15.795 2.565 ;
      RECT  14.01 2.565 14.24 2.675 ;
      RECT  15.565 2.565 15.795 3.1 ;
      RECT  15.565 3.1 16.2 3.33 ;
      RECT  10.68 1.72 11.72 1.925 ;
      RECT  10.68 1.925 12.995 1.95 ;
      RECT  11.085 1.95 12.995 2.155 ;
      RECT  11.085 2.155 11.315 3.03 ;
      RECT  12.765 2.155 12.995 3.1 ;
      RECT  10.68 3.03 11.315 3.26 ;
      RECT  12.765 3.1 13.26 3.33 ;
      RECT  7.165 1.98 10.195 2.21 ;
      RECT  9.965 2.21 10.195 2.4 ;
      RECT  7.165 2.21 7.395 2.735 ;
      RECT  9.965 2.4 10.81 2.63 ;
      RECT  9.965 2.63 10.195 3.03 ;
      RECT  9.14 3.03 10.195 3.26 ;
      RECT  16.07 2.38 20.89 2.61 ;
      RECT  16.685 2.61 16.915 3.56 ;
      RECT  12.15 1.465 13.775 1.695 ;
      RECT  13.545 1.695 13.775 3.56 ;
      RECT  12.15 3.56 16.915 3.79 ;
      RECT  8.55 2.445 9.69 2.675 ;
      RECT  8.55 2.675 8.78 3.03 ;
      RECT  5.485 1.565 6.835 1.795 ;
      RECT  6.605 1.795 6.835 3.03 ;
      RECT  5.485 1.795 5.715 3.315 ;
      RECT  6.605 3.03 8.78 3.26 ;
      RECT  1.72 3.805 4.43 4.035 ;
      RECT  4.2 4.035 4.43 4.465 ;
      RECT  4.2 4.465 6.54 4.695 ;
      RECT  4.66 4.005 7.24 4.235 ;
      RECT  11.38 4.09 15.5 4.32 ;
  END
END MDN_FDPRBQ_F_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPRBQ_1
#      Description : D-Flip Flop, pos-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPRBQ_1
  CLASS CORE ;
  FOREIGN MDN_FDPRBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 3.245 ;
      RECT  15.005 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 9.66 2.355 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  9.965 5.015 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 5.015 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  8.4 -0.14 9.52 0.14 ;
      RECT  8.845 0.14 9.075 1.005 ;
      RECT  8.44 1.005 9.48 1.235 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.6 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.465 0.37 1.85 0.6 ;
      RECT  1.465 0.6 1.695 1.005 ;
      RECT  0.18 1.005 1.695 1.235 ;
      RECT  9.965 0.37 11.93 0.6 ;
      RECT  9.965 0.6 10.195 1.465 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 0.83 ;
      RECT  1.925 0.83 6.22 1.005 ;
      RECT  1.925 1.005 7.955 1.06 ;
      RECT  5.99 1.06 7.955 1.235 ;
      RECT  1.925 1.06 2.155 1.565 ;
      RECT  7.725 1.235 7.955 1.465 ;
      RECT  7.725 1.465 10.195 1.695 ;
      RECT  1.565 1.565 2.155 1.795 ;
      RECT  1.565 1.795 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  14.94 0.37 15.29 0.6 ;
      RECT  14.94 0.6 15.17 1.005 ;
      RECT  10.68 1.005 15.17 1.235 ;
      RECT  14.445 1.235 14.675 2.125 ;
      RECT  13.885 2.125 14.675 2.355 ;
      RECT  13.885 2.355 14.115 4.02 ;
      RECT  9.105 4.02 14.115 4.25 ;
      RECT  2.42 1.29 5.0 1.52 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  12.92 1.565 13.96 1.795 ;
      RECT  11.435 1.51 11.665 1.945 ;
      RECT  9.965 1.945 11.665 2.175 ;
      RECT  9.965 2.175 10.195 3.56 ;
      RECT  3.245 1.75 4.3 1.98 ;
      RECT  3.245 1.98 3.475 3.245 ;
      RECT  3.245 3.245 5.155 3.475 ;
      RECT  4.925 3.475 5.155 3.56 ;
      RECT  4.925 3.56 13.26 3.79 ;
      RECT  7.165 2.35 7.395 3.56 ;
      RECT  5.485 1.51 5.715 2.405 ;
      RECT  3.75 2.405 5.715 2.635 ;
      RECT  5.485 2.635 5.715 3.09 ;
      RECT  5.43 3.09 5.77 3.32 ;
      RECT  12.205 1.51 12.435 2.405 ;
      RECT  10.47 2.405 12.435 2.635 ;
      RECT  12.205 2.635 12.435 3.09 ;
      RECT  12.15 3.09 12.49 3.32 ;
      RECT  2.42 3.805 4.595 4.02 ;
      RECT  2.42 4.02 6.54 4.035 ;
      RECT  4.365 4.035 6.54 4.25 ;
      RECT  6.77 4.095 8.78 4.325 ;
      RECT  6.77 4.325 7.0 4.48 ;
      RECT  4.66 4.48 7.0 4.71 ;
      RECT  11.38 4.48 13.96 4.71 ;
      RECT  7.265 4.555 10.755 4.785 ;
      RECT  7.265 4.785 7.495 5.0 ;
      RECT  10.525 4.785 10.755 5.0 ;
      RECT  0.18 4.365 4.035 4.595 ;
      RECT  1.5 4.595 1.73 5.0 ;
      RECT  3.805 4.595 4.035 5.0 ;
      RECT  1.5 5.0 1.85 5.23 ;
      RECT  3.805 5.0 7.495 5.23 ;
      RECT  10.525 5.0 13.05 5.23 ;
  END
END MDN_FDPRBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPRBQ_2
#      Description : D-Flip Flop, pos-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPRBQ_2
  CLASS CORE ;
  FOREIGN MDN_FDPRBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.16 1.565 16.2 1.795 ;
      RECT  15.565 1.795 15.795 3.245 ;
      RECT  15.16 3.245 16.2 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 9.66 2.355 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  9.965 5.015 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 5.015 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.245 4.945 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.945 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  8.4 -0.14 9.52 0.14 ;
      RECT  8.845 0.14 9.075 0.89 ;
      RECT  8.44 0.89 9.48 1.12 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.6 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  11.59 0.37 11.93 0.445 ;
      RECT  9.965 0.445 11.93 0.675 ;
      RECT  9.965 0.675 10.195 1.35 ;
      RECT  9.405 1.35 10.195 1.565 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 0.83 ;
      RECT  1.565 0.83 6.22 1.005 ;
      RECT  1.565 1.005 7.955 1.06 ;
      RECT  5.99 1.06 7.955 1.235 ;
      RECT  1.565 1.06 1.795 1.565 ;
      RECT  7.725 1.235 7.955 1.565 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  7.725 1.565 10.195 1.58 ;
      RECT  7.725 1.58 9.635 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 2.06 4.035 ;
      RECT  14.95 0.37 15.29 0.445 ;
      RECT  14.95 0.445 16.41 0.675 ;
      RECT  16.07 0.37 16.41 0.445 ;
      RECT  14.95 0.675 15.18 1.005 ;
      RECT  13.82 0.37 14.17 0.6 ;
      RECT  13.94 0.6 14.17 1.005 ;
      RECT  10.68 1.005 15.18 1.235 ;
      RECT  2.42 1.29 5.0 1.52 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  12.92 1.565 13.96 1.795 ;
      RECT  11.435 1.51 11.665 1.845 ;
      RECT  9.965 1.845 11.665 2.075 ;
      RECT  9.965 2.075 10.195 3.555 ;
      RECT  3.245 1.75 4.3 1.98 ;
      RECT  3.245 1.98 3.475 3.555 ;
      RECT  3.245 3.555 13.26 3.785 ;
      RECT  7.165 2.35 7.395 3.555 ;
      RECT  5.485 1.51 5.715 2.405 ;
      RECT  3.75 2.405 5.715 2.635 ;
      RECT  5.485 2.635 5.715 3.315 ;
      RECT  12.205 1.51 12.435 2.405 ;
      RECT  10.47 2.405 12.435 2.635 ;
      RECT  12.205 2.635 12.435 3.315 ;
      RECT  13.885 2.35 14.115 4.015 ;
      RECT  9.14 4.015 14.115 4.245 ;
      RECT  2.42 4.015 6.54 4.245 ;
      RECT  6.77 4.095 8.78 4.325 ;
      RECT  6.77 4.325 7.0 4.48 ;
      RECT  4.66 4.48 7.0 4.71 ;
      RECT  11.38 4.475 13.96 4.705 ;
      RECT  9.405 4.545 10.755 4.775 ;
      RECT  9.405 4.775 9.635 4.925 ;
      RECT  10.525 4.775 10.755 5.0 ;
      RECT  7.265 4.555 8.515 4.785 ;
      RECT  8.285 4.785 8.515 4.925 ;
      RECT  7.265 4.785 7.495 5.0 ;
      RECT  8.285 4.925 9.635 5.155 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.48 ;
      RECT  0.18 4.48 4.035 4.71 ;
      RECT  1.51 4.71 1.74 5.0 ;
      RECT  3.805 4.71 4.035 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  3.805 5.0 7.495 5.23 ;
      RECT  10.525 5.0 13.05 5.23 ;
  END
END MDN_FDPRBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPRBQ_4
#      Description : D-Flip Flop, pos-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPRBQ_4
  CLASS CORE ;
  FOREIGN MDN_FDPRBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.16 1.565 18.44 1.795 ;
      RECT  17.805 1.795 18.035 3.245 ;
      RECT  15.16 3.245 18.44 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 9.66 2.355 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  7.725 5.015 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 5.015 10.195 5.46 ;
      RECT  3.245 4.94 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.94 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  8.4 -0.14 9.52 0.14 ;
      RECT  8.845 0.14 9.075 1.005 ;
      RECT  8.44 1.005 9.48 1.235 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.6 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.675 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  11.59 0.37 11.93 0.445 ;
      RECT  9.965 0.445 11.93 0.675 ;
      RECT  9.965 0.675 10.195 1.465 ;
      RECT  9.405 1.465 10.195 1.565 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 0.83 ;
      RECT  1.565 0.83 6.22 1.005 ;
      RECT  1.565 1.005 7.955 1.06 ;
      RECT  1.565 1.06 2.06 1.235 ;
      RECT  5.99 1.06 7.955 1.235 ;
      RECT  1.565 1.235 1.795 3.805 ;
      RECT  7.725 1.235 7.955 1.565 ;
      RECT  7.725 1.565 10.195 1.695 ;
      RECT  7.725 1.695 9.635 1.795 ;
      RECT  1.565 3.805 2.06 4.035 ;
      RECT  17.19 0.37 18.65 0.6 ;
      RECT  10.68 1.005 14.675 1.235 ;
      RECT  14.445 1.235 14.675 2.405 ;
      RECT  13.885 2.405 17.53 2.635 ;
      RECT  13.885 2.635 14.115 4.005 ;
      RECT  9.14 4.005 14.115 4.235 ;
      RECT  2.42 1.29 4.945 1.52 ;
      RECT  4.715 1.52 4.945 1.85 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  12.92 1.565 13.96 1.795 ;
      RECT  11.435 1.51 11.665 1.945 ;
      RECT  9.965 1.945 11.665 2.175 ;
      RECT  9.965 2.175 10.195 3.545 ;
      RECT  3.245 1.75 4.3 1.98 ;
      RECT  3.245 1.98 3.475 3.545 ;
      RECT  3.245 3.545 13.26 3.775 ;
      RECT  7.165 2.35 7.395 3.545 ;
      RECT  5.485 1.51 5.715 2.405 ;
      RECT  3.75 2.405 5.715 2.635 ;
      RECT  5.485 2.635 5.715 3.315 ;
      RECT  12.205 1.51 12.435 2.405 ;
      RECT  10.47 2.405 12.435 2.635 ;
      RECT  12.205 2.635 12.435 3.315 ;
      RECT  2.42 4.005 6.54 4.235 ;
      RECT  6.77 4.015 8.78 4.245 ;
      RECT  6.77 4.245 7.0 4.48 ;
      RECT  4.66 4.48 7.0 4.71 ;
      RECT  11.38 4.48 13.96 4.71 ;
      RECT  7.255 4.555 10.755 4.785 ;
      RECT  7.255 4.785 7.485 5.0 ;
      RECT  10.525 4.785 10.755 5.0 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.48 ;
      RECT  0.18 4.48 4.035 4.71 ;
      RECT  1.51 4.71 1.74 5.0 ;
      RECT  3.805 4.71 4.035 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  3.805 5.0 7.485 5.23 ;
      RECT  10.525 5.0 13.05 5.23 ;
  END
END MDN_FDPRBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPRBSBQ_1
#      Description : D-Flip Flop pos-edge triggered, lo-async-clear/set, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPRBSBQ_1
  CLASS CORE ;
  FOREIGN MDN_FDPRBSBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 2.35 4.035 2.66 ;
      RECT  3.245 2.66 4.035 2.94 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.75 2.915 1.98 ;
      RECT  2.61 1.98 2.915 2.1 ;
      RECT  2.685 2.1 2.915 3.245 ;
      RECT  2.42 3.245 2.915 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 1.565 11.9 2.335 ;
      RECT  11.59 2.335 11.93 2.38 ;
      RECT  11.57 2.38 11.93 2.405 ;
      RECT  8.23 2.405 11.93 2.635 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.47 0.37 10.81 0.42 ;
      RECT  10.47 0.42 11.01 0.445 ;
      RECT  10.47 0.445 16.915 0.675 ;
      RECT  16.685 0.675 16.915 1.545 ;
      RECT  16.685 1.545 17.5 1.795 ;
      RECT  17.22 1.795 17.5 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  12.205 5.08 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.965 5.08 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 5.08 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  17.245 -0.14 18.09 0.14 ;
      RECT  17.245 0.14 17.475 1.005 ;
      RECT  17.245 1.005 17.74 1.235 ;
      RECT  9.52 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 1.005 ;
      RECT  8.44 1.005 11.72 1.235 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.52 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  9.35 0.37 9.69 0.445 ;
      RECT  7.725 0.445 9.69 0.675 ;
      RECT  7.725 0.675 7.955 1.485 ;
      RECT  6.605 1.485 7.955 1.68 ;
      RECT  5.485 1.68 7.955 1.715 ;
      RECT  5.485 1.715 6.835 1.91 ;
      RECT  5.485 1.91 5.715 3.315 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.87 0.6 5.1 0.75 ;
      RECT  1.465 0.37 2.915 0.6 ;
      RECT  2.685 0.6 2.915 0.75 ;
      RECT  1.465 0.6 1.695 1.005 ;
      RECT  2.685 0.75 5.1 0.98 ;
      RECT  0.18 1.005 1.695 1.235 ;
      RECT  5.485 0.37 6.33 0.6 ;
      RECT  5.485 0.6 5.715 1.21 ;
      RECT  1.925 1.21 5.715 1.44 ;
      RECT  1.925 1.44 2.155 1.565 ;
      RECT  1.565 1.565 2.155 1.795 ;
      RECT  1.565 1.795 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  13.62 0.93 13.96 1.005 ;
      RECT  13.62 1.005 16.2 1.235 ;
      RECT  15.86 0.93 16.2 1.005 ;
      RECT  6.2 1.005 7.24 1.235 ;
      RECT  8.845 1.565 9.48 1.795 ;
      RECT  8.845 1.795 9.075 1.945 ;
      RECT  7.165 1.945 9.075 2.175 ;
      RECT  7.165 2.175 7.395 3.03 ;
      RECT  7.165 3.03 9.48 3.26 ;
      RECT  12.205 1.565 13.265 1.795 ;
      RECT  12.205 1.795 12.435 3.24 ;
      RECT  11.085 3.235 11.315 3.24 ;
      RECT  11.085 3.24 13.26 3.47 ;
      RECT  11.085 3.47 11.315 3.56 ;
      RECT  3.805 3.56 11.315 3.79 ;
      RECT  3.805 3.79 4.035 3.805 ;
      RECT  3.245 3.805 4.035 4.035 ;
      RECT  3.245 4.035 3.475 4.365 ;
      RECT  2.74 4.365 3.475 4.595 ;
      RECT  2.74 4.595 2.97 5.0 ;
      RECT  2.63 5.0 2.97 5.23 ;
      RECT  13.885 1.565 14.735 1.795 ;
      RECT  13.885 1.795 14.115 2.4 ;
      RECT  12.71 2.4 14.115 2.63 ;
      RECT  13.885 2.63 14.115 3.24 ;
      RECT  13.885 3.24 14.73 3.47 ;
      RECT  15.16 1.565 15.795 1.795 ;
      RECT  15.565 1.795 15.795 3.7 ;
      RECT  12.205 3.7 15.795 3.93 ;
      RECT  12.205 3.93 12.435 4.025 ;
      RECT  9.14 4.025 12.435 4.255 ;
      RECT  3.955 1.67 5.0 1.9 ;
      RECT  6.27 2.27 6.505 2.66 ;
      RECT  6.27 2.66 6.91 2.94 ;
      RECT  15.005 2.35 15.235 2.66 ;
      RECT  14.37 2.66 15.235 2.94 ;
      RECT  4.66 4.02 8.78 4.25 ;
      RECT  12.92 4.16 14.675 4.39 ;
      RECT  14.445 4.39 14.675 4.925 ;
      RECT  14.445 4.925 16.41 5.155 ;
      RECT  16.07 5.155 16.41 5.23 ;
      RECT  0.18 4.365 1.74 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  15.16 4.365 17.74 4.595 ;
      RECT  3.96 4.48 6.54 4.71 ;
      RECT  7.165 4.62 14.06 4.85 ;
      RECT  7.165 4.85 7.395 5.0 ;
      RECT  13.83 4.85 14.06 5.0 ;
      RECT  4.87 5.0 7.395 5.23 ;
      RECT  13.83 5.0 14.17 5.23 ;
      LAYER METAL2 ;
      RECT  6.53 2.66 14.75 2.94 ;
      LAYER VIA12 ;
      RECT  6.59 2.67 6.85 2.93 ;
      RECT  14.43 2.67 14.69 2.93 ;
  END
END MDN_FDPRBSBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPRBSBQ_2
#      Description : D-Flip Flop pos-edge triggered, lo-async-clear/set, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPRBSBQ_2
  CLASS CORE ;
  FOREIGN MDN_FDPRBSBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.35 4.06 3.475 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.1 1.565 19.98 1.795 ;
      RECT  18.925 1.795 19.155 3.245 ;
      RECT  18.1 3.245 19.98 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 2.125 11.9 2.38 ;
      RECT  11.57 2.38 11.9 2.445 ;
      RECT  8.23 2.445 11.9 2.675 ;
      RECT  11.62 2.675 11.9 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.22 4.365 17.5 5.0 ;
      RECT  17.19 5.0 17.53 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  9.905 5.135 10.25 5.46 ;
      RECT  9.52 5.46 12.88 5.74 ;
      RECT  12.145 5.135 12.49 5.46 ;
      RECT  7.67 5.135 8.01 5.46 ;
      RECT  7.28 5.46 8.4 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  17.75 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  17.805 0.14 18.035 1.005 ;
      RECT  17.4 1.005 18.035 1.235 ;
      RECT  9.52 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 1.005 ;
      RECT  8.44 1.005 11.72 1.235 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.52 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  18.07 -0.13 18.33 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  9.35 0.37 9.69 0.445 ;
      RECT  7.725 0.445 9.69 0.675 ;
      RECT  7.725 0.675 7.955 1.465 ;
      RECT  6.605 1.465 7.955 1.675 ;
      RECT  5.485 1.675 7.955 1.695 ;
      RECT  5.485 1.695 6.835 1.905 ;
      RECT  5.485 1.905 5.715 3.53 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.87 0.6 5.1 0.75 ;
      RECT  2.63 0.37 2.97 0.445 ;
      RECT  1.565 0.445 2.97 0.675 ;
      RECT  2.74 0.675 2.97 0.75 ;
      RECT  1.565 0.675 1.795 1.565 ;
      RECT  2.74 0.75 5.1 0.98 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  5.485 0.37 6.33 0.6 ;
      RECT  5.485 0.6 5.715 1.21 ;
      RECT  2.685 1.21 5.715 1.44 ;
      RECT  2.685 1.44 2.915 1.565 ;
      RECT  2.42 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  2.42 3.245 2.915 3.475 ;
      RECT  10.47 0.37 17.53 0.6 ;
      RECT  19.43 0.37 19.77 0.6 ;
      RECT  19.43 0.6 19.66 1.005 ;
      RECT  18.31 0.37 18.65 0.6 ;
      RECT  18.42 0.6 18.65 1.005 ;
      RECT  18.42 1.005 19.66 1.235 ;
      RECT  13.035 0.83 16.92 1.06 ;
      RECT  13.035 1.06 13.265 1.565 ;
      RECT  16.69 1.06 16.92 2.405 ;
      RECT  12.205 1.565 13.265 1.795 ;
      RECT  12.205 1.795 12.435 3.245 ;
      RECT  16.07 2.405 18.65 2.635 ;
      RECT  11.38 3.245 13.26 3.475 ;
      RECT  6.2 1.005 7.24 1.235 ;
      RECT  13.62 1.29 16.2 1.52 ;
      RECT  3.96 1.67 5.0 1.9 ;
      RECT  14.39 1.75 14.73 1.98 ;
      RECT  14.445 1.98 14.675 2.415 ;
      RECT  12.71 2.415 14.675 2.645 ;
      RECT  14.445 2.645 14.675 3.525 ;
      RECT  15.005 1.75 15.5 1.98 ;
      RECT  15.005 1.98 15.235 3.755 ;
      RECT  8.285 1.565 9.48 1.795 ;
      RECT  8.285 1.795 8.515 1.94 ;
      RECT  7.165 1.94 8.515 2.17 ;
      RECT  7.165 2.17 7.395 3.1 ;
      RECT  7.165 3.1 10.195 3.33 ;
      RECT  9.965 3.33 10.195 3.755 ;
      RECT  9.965 3.755 15.235 3.985 ;
      RECT  15.565 3.245 17.74 3.475 ;
      RECT  15.565 3.475 15.795 4.365 ;
      RECT  15.16 4.365 15.795 4.595 ;
      RECT  6.045 2.345 6.275 3.56 ;
      RECT  6.045 3.56 9.635 3.79 ;
      RECT  9.405 3.79 9.635 4.215 ;
      RECT  9.405 4.215 14.675 4.445 ;
      RECT  14.445 4.445 14.675 5.0 ;
      RECT  14.445 5.0 15.29 5.23 ;
      RECT  4.66 4.02 8.78 4.25 ;
      RECT  3.96 4.48 6.54 4.71 ;
      RECT  7.165 4.675 14.06 4.905 ;
      RECT  7.165 4.905 7.395 5.0 ;
      RECT  13.83 4.905 14.06 5.0 ;
      RECT  4.87 5.0 7.395 5.23 ;
      RECT  13.83 5.0 14.17 5.23 ;
  END
END MDN_FDPRBSBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPRBSBQ_4
#      Description : D-Flip Flop pos-edge triggered, lo-async-clear/set, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPRBSBQ_4
  CLASS CORE ;
  FOREIGN MDN_FDPRBSBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.1 1.565 22.22 1.795 ;
      RECT  20.045 1.795 20.275 3.245 ;
      RECT  18.1 3.245 22.22 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 8.54 2.685 ;
      RECT  8.26 2.685 11.9 2.915 ;
      RECT  11.62 2.125 11.9 2.685 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.22 4.365 17.5 5.0 ;
      RECT  17.19 5.0 17.53 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  9.965 5.08 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 5.08 12.435 5.46 ;
      RECT  7.725 5.08 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  17.75 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.69 ;
      RECT  17.805 0.14 18.035 1.005 ;
      RECT  17.4 1.005 18.035 1.235 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 1.005 ;
      RECT  8.44 1.005 11.72 1.235 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  18.07 -0.13 18.33 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  3.8 0.37 6.33 0.6 ;
      RECT  3.8 0.6 4.03 1.005 ;
      RECT  2.475 1.005 4.03 1.235 ;
      RECT  2.475 1.235 2.705 3.53 ;
      RECT  7.725 0.37 9.69 0.6 ;
      RECT  7.725 0.6 7.955 1.0 ;
      RECT  5.485 1.0 7.955 1.23 ;
      RECT  5.485 1.23 5.715 3.53 ;
      RECT  10.47 0.37 17.53 0.6 ;
      RECT  13.035 0.83 16.915 1.06 ;
      RECT  13.035 1.06 13.265 1.565 ;
      RECT  16.685 1.06 16.915 2.405 ;
      RECT  12.205 1.565 13.265 1.795 ;
      RECT  12.205 1.795 12.435 3.24 ;
      RECT  16.07 2.405 19.775 2.635 ;
      RECT  11.38 3.24 13.265 3.47 ;
      RECT  13.62 1.29 16.2 1.52 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  14.39 1.75 14.73 1.98 ;
      RECT  14.445 1.98 14.675 2.405 ;
      RECT  12.71 2.405 14.675 2.635 ;
      RECT  14.445 2.635 14.675 3.03 ;
      RECT  14.39 3.03 14.73 3.26 ;
      RECT  14.995 1.75 15.5 1.98 ;
      RECT  14.995 1.98 15.225 3.7 ;
      RECT  7.725 1.565 9.48 1.795 ;
      RECT  7.725 1.795 7.955 2.445 ;
      RECT  7.11 2.445 7.955 2.675 ;
      RECT  7.725 2.675 7.955 3.145 ;
      RECT  7.725 3.145 10.195 3.375 ;
      RECT  9.965 3.375 10.195 3.7 ;
      RECT  9.965 3.7 15.225 3.93 ;
      RECT  20.55 2.405 21.885 2.635 ;
      RECT  4.925 2.39 5.155 3.245 ;
      RECT  3.805 3.245 5.155 3.475 ;
      RECT  3.805 3.475 4.035 3.805 ;
      RECT  2.63 0.37 2.97 0.445 ;
      RECT  1.775 0.445 2.97 0.675 ;
      RECT  1.775 0.675 2.005 3.805 ;
      RECT  1.775 3.805 4.035 4.035 ;
      RECT  6.045 2.39 6.275 3.245 ;
      RECT  6.045 3.245 7.395 3.475 ;
      RECT  6.045 3.475 6.275 3.48 ;
      RECT  7.165 3.475 7.395 3.605 ;
      RECT  7.165 3.605 9.635 3.835 ;
      RECT  9.405 3.835 9.635 4.16 ;
      RECT  9.405 4.16 14.675 4.39 ;
      RECT  14.445 4.39 14.675 5.0 ;
      RECT  14.445 5.0 15.29 5.23 ;
      RECT  15.565 3.245 17.74 3.475 ;
      RECT  15.565 3.475 15.795 4.365 ;
      RECT  15.155 4.365 15.795 4.595 ;
      RECT  4.66 4.02 6.94 4.065 ;
      RECT  4.66 4.065 8.78 4.25 ;
      RECT  6.71 4.25 8.78 4.295 ;
      RECT  3.96 4.48 6.54 4.71 ;
      RECT  7.165 4.62 14.02 4.85 ;
      RECT  7.165 4.85 7.395 5.0 ;
      RECT  13.79 4.85 14.02 5.0 ;
      RECT  4.87 5.0 7.395 5.23 ;
      RECT  13.79 5.0 14.17 5.23 ;
      RECT  19.43 5.0 20.89 5.23 ;
  END
END MDN_FDPRBSBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPSBQ_1
#      Description : D-Flip Flop pos-edge triggered, lo-async-set, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPSBQ_1
  CLASS CORE ;
  FOREIGN MDN_FDPSBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.1 5.715 2.38 ;
      RECT  4.9 2.38 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 3.245 ;
      RECT  15.005 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 1.93 13.02 2.16 ;
      RECT  8.26 2.16 8.54 2.915 ;
      RECT  12.74 2.16 13.02 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.93 12.435 5.46 ;
      RECT  12.205 5.46 15.85 5.74 ;
      RECT  14.445 4.87 14.675 5.46 ;
      RECT  7.725 5.025 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 5.025 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.0 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 1.005 ;
      RECT  12.92 1.005 14.675 1.235 ;
      RECT  8.285 -0.14 8.96 0.14 ;
      RECT  8.285 0.14 8.515 1.005 ;
      RECT  8.285 1.005 8.78 1.235 ;
      RECT  5.04 -0.14 6.16 0.14 ;
      RECT  5.43 0.14 5.77 0.465 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  9.91 0.37 10.25 0.445 ;
      RECT  9.91 0.445 14.17 0.675 ;
      RECT  13.83 0.37 14.17 0.445 ;
      RECT  7.11 0.37 7.45 0.6 ;
      RECT  7.11 0.6 7.34 0.695 ;
      RECT  3.19 0.695 7.34 0.925 ;
      RECT  9.14 1.005 11.72 1.235 ;
      RECT  2.42 1.155 6.54 1.385 ;
      RECT  6.9 1.465 11.02 1.695 ;
      RECT  7.165 1.695 7.395 2.405 ;
      RECT  6.205 2.405 7.395 2.635 ;
      RECT  7.165 2.635 7.395 3.245 ;
      RECT  6.9 3.245 9.48 3.475 ;
      RECT  13.62 1.565 14.115 1.795 ;
      RECT  13.885 1.795 14.115 3.245 ;
      RECT  11.645 2.39 11.875 3.245 ;
      RECT  11.645 3.245 14.115 3.475 ;
      RECT  13.885 3.475 14.115 4.365 ;
      RECT  13.885 4.365 15.18 4.595 ;
      RECT  14.95 4.595 15.18 5.0 ;
      RECT  14.95 5.0 15.29 5.23 ;
      RECT  3.96 1.615 5.0 1.845 ;
      RECT  10.47 2.445 10.81 2.455 ;
      RECT  9.965 2.455 10.81 2.675 ;
      RECT  9.965 2.675 10.745 2.685 ;
      RECT  9.965 2.685 10.195 3.805 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.34 ;
      RECT  1.565 2.34 2.915 2.57 ;
      RECT  1.565 2.57 1.795 3.245 ;
      RECT  2.685 2.57 2.915 3.805 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  2.685 3.805 10.195 3.835 ;
      RECT  3.805 3.605 5.71 3.805 ;
      RECT  2.685 3.835 4.035 4.035 ;
      RECT  5.48 3.835 10.195 4.035 ;
      RECT  3.96 3.145 6.54 3.375 ;
      RECT  3.245 1.615 3.475 3.53 ;
      RECT  10.68 3.805 13.26 4.035 ;
      RECT  4.365 4.095 5.0 4.325 ;
      RECT  4.365 4.325 4.595 4.365 ;
      RECT  2.42 4.365 4.595 4.595 ;
      RECT  9.91 4.365 12.995 4.595 ;
      RECT  12.765 4.595 12.995 4.995 ;
      RECT  12.765 4.995 13.975 5.0 ;
      RECT  12.765 5.0 14.17 5.225 ;
      RECT  13.83 5.225 14.17 5.23 ;
      RECT  4.925 4.565 8.515 4.795 ;
      RECT  8.285 4.795 8.515 4.995 ;
      RECT  4.925 4.795 5.155 5.0 ;
      RECT  8.285 4.995 9.54 5.0 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 1.74 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 5.155 5.23 ;
      RECT  8.285 5.0 9.69 5.225 ;
      RECT  9.35 5.225 9.69 5.23 ;
  END
END MDN_FDPSBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPSBQ_2
#      Description : D-Flip Flop pos-edge triggered, lo-async-set, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPSBQ_2
  CLASS CORE ;
  FOREIGN MDN_FDPSBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.1 5.715 2.38 ;
      RECT  4.9 2.38 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.16 1.565 16.2 1.795 ;
      RECT  15.565 1.795 15.795 3.245 ;
      RECT  15.16 3.245 16.2 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 1.925 13.02 2.155 ;
      RECT  8.26 2.155 8.54 2.915 ;
      RECT  12.74 2.155 13.02 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 5.03 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 1.005 ;
      RECT  12.92 1.005 14.675 1.235 ;
      RECT  8.285 -0.14 8.96 0.14 ;
      RECT  8.285 0.14 8.515 1.005 ;
      RECT  8.285 1.005 8.78 1.235 ;
      RECT  5.04 -0.14 6.16 0.14 ;
      RECT  5.43 0.14 5.77 0.465 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  9.91 0.375 10.25 0.445 ;
      RECT  9.91 0.445 14.17 0.675 ;
      RECT  13.83 0.37 14.17 0.445 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.14 1.005 1.74 1.235 ;
      RECT  7.11 0.37 7.45 0.6 ;
      RECT  7.11 0.6 7.34 0.695 ;
      RECT  3.19 0.695 7.34 0.925 ;
      RECT  14.95 0.37 16.41 0.6 ;
      RECT  9.14 1.005 11.72 1.235 ;
      RECT  2.42 1.155 6.54 1.385 ;
      RECT  6.9 1.465 11.02 1.695 ;
      RECT  6.9 1.695 7.13 2.405 ;
      RECT  6.215 2.405 7.13 2.635 ;
      RECT  6.9 2.635 7.13 3.245 ;
      RECT  6.9 3.245 9.48 3.475 ;
      RECT  13.62 1.565 14.115 1.795 ;
      RECT  13.885 1.795 14.115 2.405 ;
      RECT  13.885 2.405 15.075 2.635 ;
      RECT  13.885 2.635 14.115 3.245 ;
      RECT  11.59 2.445 11.93 2.675 ;
      RECT  11.645 2.675 11.875 3.245 ;
      RECT  11.645 3.245 14.115 3.475 ;
      RECT  3.96 1.615 5.0 1.845 ;
      RECT  9.965 2.44 10.81 2.67 ;
      RECT  9.965 2.67 10.195 3.805 ;
      RECT  1.72 1.695 2.915 1.925 ;
      RECT  2.685 1.925 2.915 3.805 ;
      RECT  1.72 3.805 10.195 3.88 ;
      RECT  3.805 3.65 5.72 3.805 ;
      RECT  1.72 3.88 4.035 4.035 ;
      RECT  5.49 3.88 10.195 4.035 ;
      RECT  3.96 3.145 6.54 3.375 ;
      RECT  3.245 1.645 3.475 3.53 ;
      RECT  10.68 3.805 13.26 4.035 ;
      RECT  4.365 4.11 5.055 4.34 ;
      RECT  4.365 4.34 4.595 4.365 ;
      RECT  2.42 4.365 4.595 4.595 ;
      RECT  5.485 4.36 8.515 4.57 ;
      RECT  4.925 4.57 8.515 4.59 ;
      RECT  4.925 4.59 5.715 4.8 ;
      RECT  8.285 4.59 8.515 5.0 ;
      RECT  4.925 4.8 5.155 5.0 ;
      RECT  0.18 4.365 1.74 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 5.155 5.23 ;
      RECT  8.285 5.0 9.67 5.23 ;
      RECT  11.645 4.365 12.995 4.595 ;
      RECT  11.645 4.595 11.875 4.925 ;
      RECT  12.765 4.595 12.995 5.0 ;
      RECT  9.91 4.925 11.875 5.155 ;
      RECT  12.765 5.0 14.17 5.23 ;
  END
END MDN_FDPSBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FDPSBQ_4
#      Description : D-Flip Flop pos-edge triggered, lo-async-set, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FDPSBQ_4
  CLASS CORE ;
  FOREIGN MDN_FDPSBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.1 5.715 2.38 ;
      RECT  4.9 2.38 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.16 1.565 18.44 1.795 ;
      RECT  17.805 1.795 18.035 3.245 ;
      RECT  15.16 3.245 18.44 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 1.945 13.02 2.175 ;
      RECT  8.26 2.175 8.54 2.915 ;
      RECT  12.74 2.175 13.02 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  5.485 5.075 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 5.075 7.955 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  13.27 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 1.005 ;
      RECT  12.92 1.005 14.675 1.235 ;
      RECT  8.285 -0.14 8.96 0.14 ;
      RECT  8.285 0.14 8.515 0.965 ;
      RECT  8.285 0.965 8.78 1.195 ;
      RECT  5.04 -0.14 6.16 0.14 ;
      RECT  5.43 0.14 5.77 0.465 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  13.83 0.37 14.17 0.445 ;
      RECT  9.91 0.445 14.17 0.675 ;
      RECT  17.19 0.37 17.53 0.445 ;
      RECT  17.19 0.445 18.65 0.675 ;
      RECT  18.31 0.37 18.65 0.445 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.51 0.6 1.74 1.005 ;
      RECT  0.18 1.005 1.74 1.235 ;
      RECT  7.11 0.37 7.45 0.6 ;
      RECT  7.11 0.6 7.34 0.695 ;
      RECT  3.19 0.695 7.34 0.925 ;
      RECT  9.14 0.965 11.72 1.195 ;
      RECT  2.42 1.16 6.54 1.39 ;
      RECT  6.9 1.485 11.02 1.715 ;
      RECT  7.165 1.715 7.395 2.405 ;
      RECT  6.21 2.405 7.395 2.635 ;
      RECT  7.165 2.635 7.395 3.245 ;
      RECT  6.9 3.245 9.48 3.475 ;
      RECT  13.62 1.565 14.115 1.795 ;
      RECT  13.885 1.795 14.115 2.445 ;
      RECT  13.885 2.445 17.4 2.675 ;
      RECT  13.885 2.675 14.115 3.245 ;
      RECT  11.59 2.445 11.93 2.675 ;
      RECT  11.645 2.675 11.875 3.245 ;
      RECT  11.645 3.245 14.115 3.475 ;
      RECT  3.96 1.62 5.0 1.85 ;
      RECT  9.965 2.445 10.81 2.675 ;
      RECT  9.965 2.675 10.195 3.805 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.39 ;
      RECT  1.565 2.39 2.915 2.62 ;
      RECT  1.565 2.62 1.795 3.245 ;
      RECT  2.685 2.62 2.915 3.805 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  2.685 3.805 10.195 3.835 ;
      RECT  3.805 3.605 5.715 3.805 ;
      RECT  2.685 3.835 4.035 4.035 ;
      RECT  5.485 3.835 10.195 4.035 ;
      RECT  3.96 3.145 6.54 3.375 ;
      RECT  3.245 1.62 3.475 3.53 ;
      RECT  10.68 3.805 13.26 4.035 ;
      RECT  4.365 4.065 5.005 4.295 ;
      RECT  4.365 4.295 4.595 4.365 ;
      RECT  2.42 4.365 4.595 4.595 ;
      RECT  11.645 4.365 12.995 4.595 ;
      RECT  11.645 4.595 11.875 4.925 ;
      RECT  12.765 4.595 12.995 5.0 ;
      RECT  9.91 4.925 11.875 5.155 ;
      RECT  12.765 5.0 14.17 5.23 ;
      RECT  4.925 4.615 8.515 4.845 ;
      RECT  4.925 4.845 5.155 5.0 ;
      RECT  8.285 4.845 8.515 5.0 ;
      RECT  0.17 4.365 1.74 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 5.155 5.23 ;
      RECT  8.285 5.0 9.67 5.23 ;
  END
END MDN_FDPSBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FILL1
#      Description : Filler cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FILL1
  CLASS CORE SPACER ;
  FOREIGN MDN_FILL1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.24 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.46 2.24 5.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.14 2.24 0.14 ;
    END
  END VSS
END MDN_FILL1
#-----------------------------------------------------------------------
#      Cell        : MDN_FILL16
#      Description : Filler cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FILL16
  CLASS CORE SPACER ;
  FOREIGN MDN_FILL16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 35.84 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.46 35.84 5.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.14 35.84 0.14 ;
    END
  END VSS
END MDN_FILL16
#-----------------------------------------------------------------------
#      Cell        : MDN_FILL2
#      Description : Filler cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FILL2
  CLASS CORE SPACER ;
  FOREIGN MDN_FILL2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
    END
  END VSS
END MDN_FILL2
#-----------------------------------------------------------------------
#      Cell        : MDN_FILL32
#      Description : Filler cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FILL32
  CLASS CORE SPACER ;
  FOREIGN MDN_FILL32 0 0 ;
  ORIGIN 0 0 ;
  SIZE 71.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.46 71.68 5.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.14 71.68 0.14 ;
    END
  END VSS
END MDN_FILL32
#-----------------------------------------------------------------------
#      Cell        : MDN_FILL4
#      Description : Filler cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FILL4
  CLASS CORE SPACER ;
  FOREIGN MDN_FILL4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
    END
  END VSS
END MDN_FILL4
#-----------------------------------------------------------------------
#      Cell        : MDN_FILL8
#      Description : Filler cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FILL8
  CLASS CORE SPACER ;
  FOREIGN MDN_FILL8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
    END
  END VSS
END MDN_FILL8
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL2TD1
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL2TD1
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL2TD1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.24 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.04 2.24 5.88 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.56 2.24 0.28 ;
    END
  END VSS
END MDN_RAIL2TD1
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL2TD16
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL2TD16
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL2TD16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 35.84 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.04 35.84 5.88 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.56 35.84 0.28 ;
    END
  END VSS
END MDN_RAIL2TD16
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL2TD2
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL2TD2
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL2TD2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.04 4.48 5.88 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.56 4.48 0.28 ;
    END
  END VSS
END MDN_RAIL2TD2
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL2TD32
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL2TD32
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL2TD32 0 0 ;
  ORIGIN 0 0 ;
  SIZE 71.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.04 71.68 5.88 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.56 71.68 0.28 ;
    END
  END VSS
END MDN_RAIL2TD32
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL2TD4
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL2TD4
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL2TD4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.04 8.96 5.88 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.56 8.96 0.28 ;
    END
  END VSS
END MDN_RAIL2TD4
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL2TD8
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL2TD8
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL2TD8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.04 17.92 5.88 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.56 17.92 0.28 ;
    END
  END VSS
END MDN_RAIL2TD8
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL1T1
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL1T1
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL1T1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.24 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.46 2.24 5.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.14 2.24 0.14 ;
    END
  END VSS
END MDN_RAIL1T1
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL1T16
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL1T16
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL1T16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 35.84 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.46 35.84 5.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.14 35.84 0.14 ;
    END
  END VSS
END MDN_RAIL1T16
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL1T2
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL1T2
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL1T2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
    END
  END VSS
END MDN_RAIL1T2
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL1T32
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL1T32
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL1T32 0 0 ;
  ORIGIN 0 0 ;
  SIZE 71.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.46 71.68 5.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.14 71.68 0.14 ;
    END
  END VSS
END MDN_RAIL1T32
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL1T4
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL1T4
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL1T4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
    END
  END VSS
END MDN_RAIL1T4
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL1T8
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL1T8
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL1T8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
    END
  END VSS
END MDN_RAIL1T8
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL3T1
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL3T1
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL3T1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.24 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.04 2.24 6.16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.56 2.24 0.56 ;
    END
  END VSS
END MDN_RAIL3T1
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL3T16
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL3T16
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL3T16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 35.84 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.04 35.84 6.16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.56 35.84 0.56 ;
    END
  END VSS
END MDN_RAIL3T16
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL3T2
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL3T2
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL3T2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.04 4.48 6.16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.56 4.48 0.56 ;
    END
  END VSS
END MDN_RAIL3T2
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL3T32
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL3T32
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL3T32 0 0 ;
  ORIGIN 0 0 ;
  SIZE 71.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.04 71.68 6.16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.56 71.68 0.56 ;
    END
  END VSS
END MDN_RAIL3T32
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL3T4
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL3T4
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL3T4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.04 8.96 6.16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.56 8.96 0.56 ;
    END
  END VSS
END MDN_RAIL3T4
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL3T8
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL3T8
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL3T8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.04 17.92 6.16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.56 17.92 0.56 ;
    END
  END VSS
END MDN_RAIL3T8
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL2TU1
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL2TU1
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL2TU1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.24 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.32 2.24 6.16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.28 2.24 0.56 ;
    END
  END VSS
END MDN_RAIL2TU1
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL2TU16
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL2TU16
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL2TU16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 35.84 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.32 35.84 6.16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.28 35.84 0.56 ;
    END
  END VSS
END MDN_RAIL2TU16
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL2TU2
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL2TU2
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL2TU2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.32 4.48 6.16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.28 4.48 0.56 ;
    END
  END VSS
END MDN_RAIL2TU2
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL2TU32
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL2TU32
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL2TU32 0 0 ;
  ORIGIN 0 0 ;
  SIZE 71.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.32 71.68 6.16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.28 71.68 0.56 ;
    END
  END VSS
END MDN_RAIL2TU32
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL2TU4
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL2TU4
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL2TU4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.32 8.96 6.16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.28 8.96 0.56 ;
    END
  END VSS
END MDN_RAIL2TU4
#-----------------------------------------------------------------------
#      Cell        : MDN_RAIL2TU8
#      Description : Rail cell
#      Equation    : None
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_RAIL2TU8
  CLASS CORE SPACER ;
  FOREIGN MDN_RAIL2TU8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 5.32 17.92 6.16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL2 ;
      RECT  0.0 -0.28 17.92 0.56 ;
    END
  END VSS
END MDN_RAIL2TU8
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDN_4
#      Description : D-Flip Flop w/scan, neg-edge triggered
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI)):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDN_4
  CLASS CORE ;
  FOREIGN MDN_FSDN_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 26.88 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.1 1.565 22.22 1.795 ;
      RECT  20.045 1.795 20.275 3.245 ;
      RECT  18.1 3.245 22.22 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  22.58 1.565 26.7 1.795 ;
      RECT  24.525 1.795 24.755 3.245 ;
      RECT  22.58 3.245 26.7 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.645 5.46 27.05 5.74 ;
      RECT  18.925 4.87 19.155 5.46 ;
      RECT  18.925 5.46 23.635 5.74 ;
      RECT  21.165 4.93 21.395 5.46 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  15.51 5.46 16.915 5.74 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 26.88 5.74 ;
      LAYER VIA12 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  20.31 5.47 20.57 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  22.55 5.47 22.81 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 27.05 0.14 ;
      RECT  21.165 0.14 21.395 0.73 ;
      RECT  23.405 0.14 23.635 0.73 ;
      RECT  25.645 0.14 25.875 0.73 ;
      RECT  17.75 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  15.51 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  5.485 -0.14 6.89 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.24 -0.14 2.915 0.14 ;
      RECT  2.685 0.14 2.915 1.005 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 26.88 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  22.55 -0.13 22.81 0.13 ;
      RECT  23.11 -0.13 23.37 0.13 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  24.79 -0.13 25.05 0.13 ;
      RECT  25.35 -0.13 25.61 0.13 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  18.07 -0.13 18.33 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  12.765 0.37 15.295 0.6 ;
      RECT  12.765 0.6 12.995 1.005 ;
      RECT  12.205 1.005 12.995 1.235 ;
      RECT  12.205 1.235 12.435 1.565 ;
      RECT  9.965 1.565 12.435 1.795 ;
      RECT  9.965 1.795 10.195 2.34 ;
      RECT  9.35 2.34 10.195 2.57 ;
      RECT  16.07 0.37 16.41 0.6 ;
      RECT  16.07 0.6 16.3 1.005 ;
      RECT  14.39 1.005 16.3 1.235 ;
      RECT  26.15 0.37 26.49 0.6 ;
      RECT  26.15 0.6 26.38 1.01 ;
      RECT  23.91 0.37 25.37 0.6 ;
      RECT  23.91 0.6 24.14 1.005 ;
      RECT  25.14 0.6 25.37 1.01 ;
      RECT  22.79 0.37 23.13 0.6 ;
      RECT  22.9 0.6 23.13 1.005 ;
      RECT  17.245 1.005 24.14 1.235 ;
      RECT  25.14 1.01 26.38 1.24 ;
      RECT  17.245 1.235 17.475 3.24 ;
      RECT  17.245 3.24 17.74 3.47 ;
      RECT  7.01 0.445 9.635 0.675 ;
      RECT  7.01 0.675 7.24 0.89 ;
      RECT  9.405 0.675 9.635 1.005 ;
      RECT  6.9 0.89 7.24 1.12 ;
      RECT  9.405 1.005 11.72 1.235 ;
      RECT  7.685 1.005 8.78 1.01 ;
      RECT  7.68 1.01 8.78 1.015 ;
      RECT  7.675 1.015 8.78 1.02 ;
      RECT  7.67 1.02 8.78 1.025 ;
      RECT  7.665 1.025 8.78 1.03 ;
      RECT  7.66 1.03 8.78 1.035 ;
      RECT  7.655 1.035 8.78 1.04 ;
      RECT  7.65 1.04 8.78 1.045 ;
      RECT  7.645 1.045 8.78 1.05 ;
      RECT  7.64 1.05 8.78 1.055 ;
      RECT  7.635 1.055 8.78 1.06 ;
      RECT  7.63 1.06 8.78 1.065 ;
      RECT  7.625 1.065 8.78 1.07 ;
      RECT  7.62 1.07 8.78 1.075 ;
      RECT  7.615 1.075 8.78 1.08 ;
      RECT  7.61 1.08 8.78 1.085 ;
      RECT  7.605 1.085 8.78 1.09 ;
      RECT  7.6 1.09 8.78 1.095 ;
      RECT  7.595 1.095 8.78 1.1 ;
      RECT  7.59 1.1 8.78 1.105 ;
      RECT  7.585 1.105 8.78 1.11 ;
      RECT  7.58 1.11 8.78 1.115 ;
      RECT  7.575 1.115 8.78 1.12 ;
      RECT  7.57 1.12 8.78 1.125 ;
      RECT  7.565 1.125 8.78 1.13 ;
      RECT  7.56 1.13 8.78 1.135 ;
      RECT  7.555 1.135 8.78 1.14 ;
      RECT  7.55 1.14 8.78 1.145 ;
      RECT  7.545 1.145 8.78 1.15 ;
      RECT  7.54 1.15 8.78 1.155 ;
      RECT  7.535 1.155 8.78 1.16 ;
      RECT  7.53 1.16 8.78 1.165 ;
      RECT  7.525 1.165 8.78 1.17 ;
      RECT  7.52 1.17 8.78 1.175 ;
      RECT  7.515 1.175 8.78 1.18 ;
      RECT  7.51 1.18 8.78 1.185 ;
      RECT  7.505 1.185 8.78 1.19 ;
      RECT  7.5 1.19 8.78 1.195 ;
      RECT  7.495 1.195 8.78 1.2 ;
      RECT  7.49 1.2 8.78 1.205 ;
      RECT  7.485 1.205 8.78 1.21 ;
      RECT  7.48 1.21 8.78 1.215 ;
      RECT  7.475 1.215 8.78 1.22 ;
      RECT  7.47 1.22 8.78 1.225 ;
      RECT  7.465 1.225 8.78 1.23 ;
      RECT  7.46 1.23 8.78 1.235 ;
      RECT  7.455 1.235 7.78 1.24 ;
      RECT  7.45 1.24 7.775 1.245 ;
      RECT  7.445 1.245 7.77 1.25 ;
      RECT  7.44 1.25 7.765 1.255 ;
      RECT  7.435 1.255 7.76 1.26 ;
      RECT  7.43 1.26 7.755 1.265 ;
      RECT  7.425 1.265 7.75 1.27 ;
      RECT  7.42 1.27 7.745 1.275 ;
      RECT  7.415 1.275 7.74 1.28 ;
      RECT  7.41 1.28 7.735 1.285 ;
      RECT  7.405 1.285 7.73 1.29 ;
      RECT  7.4 1.29 7.725 1.295 ;
      RECT  7.395 1.295 7.72 1.3 ;
      RECT  7.39 1.3 7.715 1.305 ;
      RECT  7.385 1.305 7.71 1.31 ;
      RECT  7.38 1.31 7.705 1.315 ;
      RECT  7.375 1.315 7.7 1.32 ;
      RECT  7.37 1.32 7.695 1.325 ;
      RECT  7.365 1.325 7.69 1.33 ;
      RECT  7.36 1.33 7.685 1.335 ;
      RECT  7.355 1.335 7.68 1.34 ;
      RECT  7.35 1.34 7.675 1.345 ;
      RECT  7.345 1.345 7.67 1.35 ;
      RECT  7.34 1.35 7.665 1.355 ;
      RECT  7.335 1.355 7.66 1.36 ;
      RECT  7.33 1.36 7.655 1.365 ;
      RECT  7.325 1.365 7.65 1.37 ;
      RECT  7.32 1.37 7.645 1.375 ;
      RECT  3.245 1.005 6.46 1.01 ;
      RECT  3.245 1.01 6.465 1.015 ;
      RECT  3.245 1.015 6.47 1.02 ;
      RECT  3.245 1.02 6.475 1.025 ;
      RECT  3.245 1.025 6.48 1.03 ;
      RECT  3.245 1.03 6.485 1.035 ;
      RECT  3.245 1.035 6.49 1.04 ;
      RECT  3.245 1.04 6.495 1.045 ;
      RECT  3.245 1.045 6.5 1.05 ;
      RECT  3.245 1.05 6.505 1.055 ;
      RECT  3.245 1.055 6.51 1.06 ;
      RECT  3.245 1.06 6.515 1.065 ;
      RECT  3.245 1.065 6.52 1.07 ;
      RECT  3.245 1.07 6.525 1.075 ;
      RECT  3.245 1.075 6.53 1.08 ;
      RECT  3.245 1.08 6.535 1.085 ;
      RECT  3.245 1.085 6.54 1.09 ;
      RECT  3.245 1.09 6.545 1.095 ;
      RECT  3.245 1.095 6.55 1.1 ;
      RECT  3.245 1.1 6.555 1.105 ;
      RECT  3.245 1.105 6.56 1.11 ;
      RECT  3.245 1.11 6.565 1.115 ;
      RECT  3.245 1.115 6.57 1.12 ;
      RECT  3.245 1.12 6.575 1.125 ;
      RECT  3.245 1.125 6.58 1.13 ;
      RECT  3.245 1.13 6.585 1.135 ;
      RECT  3.245 1.135 6.59 1.14 ;
      RECT  3.245 1.14 6.595 1.145 ;
      RECT  3.245 1.145 6.6 1.15 ;
      RECT  3.245 1.15 6.605 1.155 ;
      RECT  3.245 1.155 6.61 1.16 ;
      RECT  3.245 1.16 6.615 1.165 ;
      RECT  3.245 1.165 6.62 1.17 ;
      RECT  3.245 1.17 6.625 1.175 ;
      RECT  3.245 1.175 6.63 1.18 ;
      RECT  3.245 1.18 6.635 1.185 ;
      RECT  3.245 1.185 6.64 1.19 ;
      RECT  3.245 1.19 6.645 1.195 ;
      RECT  3.245 1.195 6.65 1.2 ;
      RECT  3.245 1.2 6.655 1.205 ;
      RECT  3.245 1.205 6.66 1.21 ;
      RECT  3.245 1.21 6.665 1.215 ;
      RECT  3.245 1.215 6.67 1.22 ;
      RECT  3.245 1.22 6.675 1.225 ;
      RECT  3.245 1.225 6.68 1.23 ;
      RECT  3.245 1.23 6.685 1.235 ;
      RECT  6.355 1.235 6.69 1.24 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  6.36 1.24 6.695 1.245 ;
      RECT  6.365 1.245 6.7 1.25 ;
      RECT  6.37 1.25 6.705 1.255 ;
      RECT  6.375 1.255 6.71 1.26 ;
      RECT  6.38 1.26 6.715 1.265 ;
      RECT  6.385 1.265 6.72 1.27 ;
      RECT  6.39 1.27 6.725 1.275 ;
      RECT  6.395 1.275 6.73 1.28 ;
      RECT  6.4 1.28 6.735 1.285 ;
      RECT  6.405 1.285 6.74 1.29 ;
      RECT  6.41 1.29 6.745 1.295 ;
      RECT  6.415 1.295 6.75 1.3 ;
      RECT  6.42 1.3 6.755 1.305 ;
      RECT  6.425 1.305 6.76 1.31 ;
      RECT  6.43 1.31 6.765 1.315 ;
      RECT  6.435 1.315 6.77 1.32 ;
      RECT  6.44 1.32 6.775 1.325 ;
      RECT  6.445 1.325 6.78 1.33 ;
      RECT  6.45 1.33 6.785 1.335 ;
      RECT  6.455 1.335 6.79 1.34 ;
      RECT  6.46 1.34 6.795 1.345 ;
      RECT  6.465 1.345 6.8 1.35 ;
      RECT  6.47 1.35 6.805 1.355 ;
      RECT  6.475 1.355 6.81 1.36 ;
      RECT  6.48 1.36 6.815 1.365 ;
      RECT  6.485 1.365 6.82 1.37 ;
      RECT  6.49 1.37 6.825 1.375 ;
      RECT  6.495 1.375 7.64 1.38 ;
      RECT  6.5 1.38 7.635 1.385 ;
      RECT  6.505 1.385 7.63 1.39 ;
      RECT  6.51 1.39 7.625 1.395 ;
      RECT  6.515 1.395 7.62 1.4 ;
      RECT  6.52 1.4 7.615 1.405 ;
      RECT  6.525 1.405 7.61 1.41 ;
      RECT  6.53 1.41 7.605 1.415 ;
      RECT  6.535 1.415 7.6 1.42 ;
      RECT  6.54 1.42 7.595 1.425 ;
      RECT  6.545 1.425 7.59 1.43 ;
      RECT  6.55 1.43 7.585 1.435 ;
      RECT  6.555 1.435 7.58 1.44 ;
      RECT  6.56 1.44 7.575 1.445 ;
      RECT  6.565 1.445 7.57 1.45 ;
      RECT  6.57 1.45 7.565 1.455 ;
      RECT  6.575 1.455 7.56 1.46 ;
      RECT  6.58 1.46 7.555 1.465 ;
      RECT  6.585 1.465 7.55 1.47 ;
      RECT  6.59 1.47 7.545 1.475 ;
      RECT  6.595 1.475 7.54 1.48 ;
      RECT  6.6 1.48 7.535 1.485 ;
      RECT  6.605 1.485 7.53 1.49 ;
      RECT  6.61 1.49 7.525 1.495 ;
      RECT  6.615 1.495 7.52 1.5 ;
      RECT  6.62 1.5 7.515 1.505 ;
      RECT  6.625 1.505 7.51 1.51 ;
      RECT  6.63 1.51 7.505 1.515 ;
      RECT  6.635 1.515 7.5 1.52 ;
      RECT  6.64 1.52 7.495 1.525 ;
      RECT  6.645 1.525 7.49 1.53 ;
      RECT  6.65 1.53 7.485 1.535 ;
      RECT  6.655 1.535 7.48 1.54 ;
      RECT  6.66 1.54 7.475 1.545 ;
      RECT  6.665 1.545 7.47 1.55 ;
      RECT  6.67 1.55 7.465 1.555 ;
      RECT  6.675 1.555 7.46 1.56 ;
      RECT  6.68 1.56 7.455 1.565 ;
      RECT  1.72 1.565 3.475 1.795 ;
      RECT  6.685 1.565 7.45 1.57 ;
      RECT  6.69 1.57 7.445 1.575 ;
      RECT  6.695 1.575 7.44 1.58 ;
      RECT  6.7 1.58 7.435 1.585 ;
      RECT  6.705 1.585 7.43 1.59 ;
      RECT  6.71 1.59 7.425 1.595 ;
      RECT  6.715 1.595 7.42 1.6 ;
      RECT  6.72 1.6 7.415 1.605 ;
      RECT  4.66 1.565 5.15 1.795 ;
      RECT  4.92 1.795 5.15 3.245 ;
      RECT  2.685 2.35 2.915 3.245 ;
      RECT  2.685 3.245 5.15 3.475 ;
      RECT  12.92 1.565 13.96 1.795 ;
      RECT  14.445 1.565 15.5 1.795 ;
      RECT  14.445 1.795 14.675 3.245 ;
      RECT  12.195 3.245 14.675 3.475 ;
      RECT  12.195 3.475 12.425 3.78 ;
      RECT  12.045 3.78 12.425 4.06 ;
      RECT  12.195 4.06 12.425 4.365 ;
      RECT  11.705 4.365 12.425 4.595 ;
      RECT  11.705 4.595 11.935 5.0 ;
      RECT  11.59 5.0 11.935 5.23 ;
      RECT  5.485 1.75 6.54 1.98 ;
      RECT  5.485 1.98 5.715 3.245 ;
      RECT  5.485 3.245 7.39 3.475 ;
      RECT  7.16 3.475 7.39 3.78 ;
      RECT  7.16 3.78 8.12 4.06 ;
      RECT  7.725 1.695 7.955 2.405 ;
      RECT  5.99 2.405 7.955 2.635 ;
      RECT  7.725 2.635 7.955 3.53 ;
      RECT  11.635 2.335 14.17 2.565 ;
      RECT  11.635 2.565 11.865 3.245 ;
      RECT  8.285 1.565 9.48 1.795 ;
      RECT  8.285 1.795 8.515 3.245 ;
      RECT  8.285 3.245 11.865 3.475 ;
      RECT  1.005 3.805 2.76 4.035 ;
      RECT  1.005 4.035 1.235 4.365 ;
      RECT  0.18 4.365 1.235 4.595 ;
      RECT  3.19 3.805 6.835 4.035 ;
      RECT  6.605 4.035 6.835 4.365 ;
      RECT  6.605 4.365 7.245 4.595 ;
      RECT  8.44 3.805 11.72 4.035 ;
      RECT  12.92 3.805 15.5 4.035 ;
      RECT  20.66 4.36 21.855 4.59 ;
      RECT  20.66 4.59 20.89 5.0 ;
      RECT  21.625 4.59 21.855 5.0 ;
      RECT  18.42 4.36 19.62 4.59 ;
      RECT  18.42 4.59 18.65 5.0 ;
      RECT  19.39 4.59 19.62 5.0 ;
      RECT  15.86 1.565 16.35 1.795 ;
      RECT  16.12 1.795 16.35 4.365 ;
      RECT  13.335 4.365 17.42 4.595 ;
      RECT  13.335 4.595 13.565 5.0 ;
      RECT  17.19 4.595 17.42 5.0 ;
      RECT  12.71 5.0 13.565 5.23 ;
      RECT  17.19 5.0 18.65 5.23 ;
      RECT  19.39 5.0 20.89 5.23 ;
      RECT  21.625 5.0 21.98 5.23 ;
      RECT  1.72 4.365 4.3 4.595 ;
      RECT  9.46 4.365 11.02 4.595 ;
      RECT  9.46 4.595 9.69 5.0 ;
      RECT  7.11 5.0 9.69 5.23 ;
      RECT  1.51 5.0 5.21 5.23 ;
      RECT  14.39 5.0 16.41 5.23 ;
      LAYER METAL2 ;
      RECT  7.74 3.78 12.425 4.06 ;
      LAYER VIA12 ;
      RECT  7.8 3.79 8.06 4.05 ;
      RECT  12.105 3.79 12.365 4.05 ;
  END
END MDN_FSDN_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDN_1
#      Description : D-Flip Flop w/scan, neg-edge triggered
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI)):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDN_1
  CLASS CORE ;
  FOREIGN MDN_FSDN_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.1 1.565 18.595 1.795 ;
      RECT  18.365 1.795 18.595 3.245 ;
      RECT  18.1 3.245 18.595 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.245 1.565 17.74 1.795 ;
      RECT  17.245 1.795 17.475 3.245 ;
      RECT  17.245 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.24 5.46 17.36 5.74 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.24 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  5.485 -0.14 6.89 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.07 -0.14 2.915 0.14 ;
      RECT  2.685 0.14 2.915 1.005 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  14.95 0.37 15.29 0.45 ;
      RECT  12.765 0.45 15.29 0.68 ;
      RECT  12.765 0.68 12.995 1.005 ;
      RECT  12.205 1.005 12.995 1.235 ;
      RECT  12.205 1.235 12.435 1.565 ;
      RECT  9.35 0.37 9.69 0.6 ;
      RECT  9.46 0.6 9.69 1.005 ;
      RECT  9.46 1.005 10.755 1.235 ;
      RECT  10.525 1.235 10.755 1.565 ;
      RECT  10.525 1.565 12.435 1.795 ;
      RECT  17.19 0.37 17.53 0.6 ;
      RECT  17.19 0.6 17.42 1.005 ;
      RECT  16.07 0.37 16.41 0.6 ;
      RECT  16.18 0.6 16.41 1.005 ;
      RECT  14.39 1.005 17.42 1.235 ;
      RECT  6.045 0.445 8.67 0.675 ;
      RECT  6.045 0.675 6.275 1.005 ;
      RECT  8.44 0.675 8.67 1.005 ;
      RECT  3.245 1.005 6.275 1.235 ;
      RECT  8.44 1.005 8.78 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  1.72 1.565 3.475 1.795 ;
      RECT  6.9 0.98 8.21 1.26 ;
      RECT  10.985 0.98 11.72 1.26 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 3.245 ;
      RECT  2.685 2.35 2.915 3.245 ;
      RECT  2.685 3.245 5.155 3.475 ;
      RECT  5.485 1.565 6.54 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  5.485 3.245 7.47 3.475 ;
      RECT  7.09 3.22 7.47 3.245 ;
      RECT  7.09 3.475 7.47 3.5 ;
      RECT  12.92 1.565 13.96 1.795 ;
      RECT  14.445 1.565 15.5 1.795 ;
      RECT  14.445 1.795 14.675 3.245 ;
      RECT  12.13 3.22 12.51 3.245 ;
      RECT  12.13 3.245 14.675 3.475 ;
      RECT  12.13 3.475 12.51 3.5 ;
      RECT  12.205 3.5 12.435 4.365 ;
      RECT  11.7 4.365 12.435 4.595 ;
      RECT  11.7 4.595 11.93 5.0 ;
      RECT  11.59 5.0 11.93 5.23 ;
      RECT  15.86 1.565 16.355 1.795 ;
      RECT  16.125 1.795 16.355 4.365 ;
      RECT  13.325 4.365 17.475 4.595 ;
      RECT  13.325 4.595 13.555 5.0 ;
      RECT  17.245 4.595 17.475 5.0 ;
      RECT  12.71 5.0 13.555 5.23 ;
      RECT  17.245 5.0 18.65 5.23 ;
      RECT  7.725 1.51 7.955 2.125 ;
      RECT  6.045 2.125 7.955 2.355 ;
      RECT  6.045 2.355 6.275 2.68 ;
      RECT  7.725 2.355 7.955 3.53 ;
      RECT  13.885 2.365 14.115 2.685 ;
      RECT  11.645 2.685 14.115 2.915 ;
      RECT  11.645 2.915 11.875 3.245 ;
      RECT  8.285 1.565 9.48 1.795 ;
      RECT  8.285 1.795 8.515 3.245 ;
      RECT  8.285 3.245 11.875 3.475 ;
      RECT  1.005 3.805 2.76 4.035 ;
      RECT  1.005 4.035 1.235 4.365 ;
      RECT  0.18 4.365 1.235 4.595 ;
      RECT  3.19 3.805 6.835 4.035 ;
      RECT  6.605 4.035 6.835 4.365 ;
      RECT  6.605 4.365 7.24 4.595 ;
      RECT  8.44 3.805 11.72 4.035 ;
      RECT  12.92 3.805 15.57 4.035 ;
      RECT  1.72 4.365 4.3 4.595 ;
      RECT  9.46 4.365 11.02 4.595 ;
      RECT  9.46 4.595 9.69 5.0 ;
      RECT  7.11 5.0 9.69 5.23 ;
      RECT  1.51 5.0 5.21 5.23 ;
      RECT  14.39 5.0 16.41 5.23 ;
      LAYER METAL2 ;
      RECT  7.83 0.98 11.39 1.26 ;
      RECT  7.09 3.22 12.51 3.5 ;
      LAYER VIA12 ;
      RECT  7.89 0.99 8.15 1.25 ;
      RECT  11.07 0.99 11.33 1.25 ;
      RECT  7.15 3.23 7.41 3.49 ;
      RECT  12.19 3.23 12.45 3.49 ;
  END
END MDN_FSDN_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDN_2
#      Description : D-Flip Flop w/scan, neg-edge triggered
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI)):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDN_2
  CLASS CORE ;
  FOREIGN MDN_FSDN_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.64 1.565 20.68 1.795 ;
      RECT  20.045 1.795 20.275 3.245 ;
      RECT  19.64 3.245 20.68 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.4 1.565 18.44 1.795 ;
      RECT  17.805 1.795 18.035 3.245 ;
      RECT  17.4 3.245 18.44 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.87 19.155 5.46 ;
      RECT  18.925 5.46 22.57 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  15.51 5.46 16.915 5.74 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  20.31 5.47 20.57 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  16.24 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  5.485 -0.14 6.89 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.07 -0.14 2.915 0.14 ;
      RECT  2.685 0.14 2.915 1.005 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  18.07 -0.13 18.33 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  14.95 0.37 15.29 0.445 ;
      RECT  12.765 0.445 15.29 0.675 ;
      RECT  12.765 0.675 12.995 1.005 ;
      RECT  12.205 1.005 12.995 1.235 ;
      RECT  12.205 1.235 12.435 1.565 ;
      RECT  9.35 0.37 9.69 0.6 ;
      RECT  9.46 0.6 9.69 1.005 ;
      RECT  9.46 1.005 10.755 1.235 ;
      RECT  10.525 1.235 10.755 1.565 ;
      RECT  10.525 1.565 12.435 1.795 ;
      RECT  17.19 0.37 18.65 0.6 ;
      RECT  17.19 0.6 17.42 1.005 ;
      RECT  16.07 0.37 16.41 0.6 ;
      RECT  16.18 0.6 16.41 1.005 ;
      RECT  14.39 1.005 17.42 1.235 ;
      RECT  6.045 0.445 8.515 0.675 ;
      RECT  6.045 0.675 6.275 1.005 ;
      RECT  8.285 0.675 8.515 1.005 ;
      RECT  3.245 1.005 6.275 1.235 ;
      RECT  8.285 1.005 8.78 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  1.72 1.565 3.475 1.795 ;
      RECT  7.675 0.98 8.055 1.005 ;
      RECT  6.86 1.005 8.055 1.235 ;
      RECT  7.675 1.235 8.055 1.26 ;
      RECT  10.995 0.98 11.715 1.005 ;
      RECT  10.995 1.005 11.72 1.235 ;
      RECT  10.995 1.235 11.715 1.26 ;
      RECT  12.92 1.56 13.955 1.565 ;
      RECT  12.92 1.565 13.96 1.795 ;
      RECT  12.92 1.795 13.955 1.8 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 3.245 ;
      RECT  2.685 2.35 2.915 3.245 ;
      RECT  2.685 3.245 5.155 3.475 ;
      RECT  5.485 1.565 6.54 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  5.485 3.245 7.395 3.475 ;
      RECT  7.165 3.475 7.395 3.805 ;
      RECT  7.165 3.805 8.21 4.035 ;
      RECT  7.83 3.78 8.21 3.805 ;
      RECT  7.83 4.035 8.21 4.06 ;
      RECT  14.445 1.565 15.5 1.795 ;
      RECT  14.445 1.795 14.675 3.245 ;
      RECT  12.205 3.245 14.675 3.475 ;
      RECT  12.205 3.475 12.435 3.78 ;
      RECT  12.055 3.78 12.435 4.06 ;
      RECT  12.205 4.06 12.435 4.365 ;
      RECT  11.59 4.365 12.435 4.595 ;
      RECT  11.59 4.595 11.82 5.0 ;
      RECT  11.59 5.0 11.93 5.23 ;
      RECT  15.86 1.565 16.355 1.795 ;
      RECT  16.125 1.795 16.355 4.365 ;
      RECT  13.325 4.365 19.66 4.595 ;
      RECT  13.325 4.595 13.555 4.925 ;
      RECT  19.43 4.595 19.66 5.0 ;
      RECT  12.71 4.925 13.555 5.155 ;
      RECT  19.43 5.0 20.89 5.23 ;
      RECT  12.71 5.155 13.05 5.23 ;
      RECT  7.725 1.51 7.955 2.125 ;
      RECT  6.045 2.125 7.955 2.355 ;
      RECT  6.045 2.355 6.275 2.69 ;
      RECT  7.725 2.355 7.955 3.53 ;
      RECT  13.885 2.36 14.115 2.685 ;
      RECT  11.645 2.685 14.115 2.915 ;
      RECT  11.645 2.915 11.875 3.245 ;
      RECT  8.285 1.565 9.48 1.795 ;
      RECT  8.285 1.795 8.515 3.245 ;
      RECT  8.285 3.245 11.875 3.475 ;
      RECT  1.005 3.805 2.76 4.035 ;
      RECT  1.005 4.035 1.235 4.365 ;
      RECT  0.18 4.365 1.235 4.595 ;
      RECT  3.19 3.805 6.835 4.035 ;
      RECT  6.605 4.035 6.835 4.365 ;
      RECT  6.605 4.365 7.24 4.595 ;
      RECT  8.44 3.805 11.72 4.035 ;
      RECT  12.92 3.805 15.5 4.035 ;
      RECT  1.72 4.365 4.3 4.595 ;
      RECT  9.46 4.365 11.02 4.595 ;
      RECT  9.46 4.595 9.69 4.925 ;
      RECT  7.11 4.925 9.69 5.155 ;
      RECT  7.11 5.155 7.45 5.23 ;
      RECT  9.35 5.155 9.69 5.23 ;
      RECT  1.51 4.925 5.21 5.155 ;
      RECT  1.51 5.155 1.85 5.23 ;
      RECT  4.87 5.155 5.21 5.23 ;
      RECT  14.39 4.925 16.41 5.155 ;
      RECT  16.07 5.155 16.41 5.23 ;
      LAYER METAL2 ;
      RECT  7.675 0.98 11.39 1.26 ;
      RECT  7.83 3.78 12.435 4.06 ;
      LAYER VIA12 ;
      RECT  7.735 0.99 7.995 1.25 ;
      RECT  11.07 0.99 11.33 1.25 ;
      RECT  7.89 3.79 8.15 4.05 ;
      RECT  12.115 3.79 12.375 4.05 ;
  END
END MDN_FSDN_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNQ_1
#      Description : D-Flip Flop w/scan, neg-edge triggered, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNQ_1
  CLASS CORE ;
  FOREIGN MDN_FSDNQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.98 2.35 15.26 3.475 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.245 1.565 17.74 1.795 ;
      RECT  17.245 1.795 17.475 3.245 ;
      RECT  17.245 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.94 14.675 5.46 ;
      RECT  14.445 5.46 18.09 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  5.485 4.93 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 18.09 0.14 ;
      RECT  14.445 0.14 14.675 0.6 ;
      RECT  16.685 0.14 16.915 0.6 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.605 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 4.3 1.12 ;
      RECT  3.245 0.89 4.3 1.005 ;
      RECT  0.18 1.12 3.475 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 5.21 0.6 ;
      RECT  5.99 0.37 7.955 0.6 ;
      RECT  7.725 0.6 7.955 3.055 ;
      RECT  7.67 3.055 8.01 3.285 ;
      RECT  10.525 0.37 14.17 0.6 ;
      RECT  10.525 0.6 10.755 0.835 ;
      RECT  8.23 0.37 8.57 0.6 ;
      RECT  8.34 0.6 8.57 0.835 ;
      RECT  8.34 0.835 10.755 1.065 ;
      RECT  17.19 0.37 17.53 0.6 ;
      RECT  17.19 0.6 17.42 0.83 ;
      RECT  16.07 0.37 16.41 0.6 ;
      RECT  16.18 0.6 16.41 0.83 ;
      RECT  11.085 0.83 17.42 1.06 ;
      RECT  11.085 1.06 11.315 1.295 ;
      RECT  10.525 1.295 11.315 1.525 ;
      RECT  10.525 1.525 10.755 3.03 ;
      RECT  10.525 3.03 11.02 3.26 ;
      RECT  4.745 1.005 7.24 1.01 ;
      RECT  4.74 1.01 7.24 1.015 ;
      RECT  4.735 1.015 7.24 1.02 ;
      RECT  4.73 1.02 7.24 1.025 ;
      RECT  4.725 1.025 7.24 1.03 ;
      RECT  4.72 1.03 7.24 1.035 ;
      RECT  4.715 1.035 7.24 1.04 ;
      RECT  4.71 1.04 7.24 1.045 ;
      RECT  4.705 1.045 7.24 1.05 ;
      RECT  4.7 1.05 7.24 1.055 ;
      RECT  4.695 1.055 7.24 1.06 ;
      RECT  4.69 1.06 7.24 1.065 ;
      RECT  4.685 1.065 7.24 1.07 ;
      RECT  4.68 1.07 7.24 1.075 ;
      RECT  4.675 1.075 7.24 1.08 ;
      RECT  4.67 1.08 7.24 1.085 ;
      RECT  4.665 1.085 7.24 1.09 ;
      RECT  4.66 1.09 7.24 1.095 ;
      RECT  4.655 1.095 7.24 1.1 ;
      RECT  4.65 1.1 7.24 1.105 ;
      RECT  4.645 1.105 7.24 1.11 ;
      RECT  4.64 1.11 7.24 1.115 ;
      RECT  4.635 1.115 7.24 1.12 ;
      RECT  4.63 1.12 7.24 1.125 ;
      RECT  4.625 1.125 7.24 1.13 ;
      RECT  4.62 1.13 7.24 1.135 ;
      RECT  4.615 1.135 7.24 1.14 ;
      RECT  4.61 1.14 7.24 1.145 ;
      RECT  4.605 1.145 7.24 1.15 ;
      RECT  4.6 1.15 7.24 1.155 ;
      RECT  4.595 1.155 7.24 1.16 ;
      RECT  4.59 1.16 7.24 1.165 ;
      RECT  4.585 1.165 7.24 1.17 ;
      RECT  4.58 1.17 7.24 1.175 ;
      RECT  4.575 1.175 7.24 1.18 ;
      RECT  4.57 1.18 7.24 1.185 ;
      RECT  4.565 1.185 7.24 1.19 ;
      RECT  4.56 1.19 7.24 1.195 ;
      RECT  4.555 1.195 7.24 1.2 ;
      RECT  4.55 1.2 7.24 1.205 ;
      RECT  4.545 1.205 7.24 1.21 ;
      RECT  4.54 1.21 7.24 1.215 ;
      RECT  4.535 1.215 7.24 1.22 ;
      RECT  4.53 1.22 7.24 1.225 ;
      RECT  4.525 1.225 7.24 1.23 ;
      RECT  4.52 1.23 7.24 1.235 ;
      RECT  4.515 1.235 4.84 1.24 ;
      RECT  4.51 1.24 4.835 1.245 ;
      RECT  4.505 1.245 4.83 1.25 ;
      RECT  4.5 1.25 4.825 1.255 ;
      RECT  4.495 1.255 4.82 1.26 ;
      RECT  4.49 1.26 4.815 1.265 ;
      RECT  4.485 1.265 4.81 1.27 ;
      RECT  4.48 1.27 4.805 1.275 ;
      RECT  4.475 1.275 4.8 1.28 ;
      RECT  4.47 1.28 4.795 1.285 ;
      RECT  4.465 1.285 4.79 1.29 ;
      RECT  4.46 1.29 4.785 1.295 ;
      RECT  4.455 1.295 4.78 1.3 ;
      RECT  4.45 1.3 4.775 1.305 ;
      RECT  4.445 1.305 4.77 1.31 ;
      RECT  4.44 1.31 4.765 1.315 ;
      RECT  4.435 1.315 4.76 1.32 ;
      RECT  4.43 1.32 4.755 1.325 ;
      RECT  4.425 1.325 4.75 1.33 ;
      RECT  4.42 1.33 4.745 1.335 ;
      RECT  4.415 1.335 4.74 1.34 ;
      RECT  4.41 1.34 4.735 1.345 ;
      RECT  4.405 1.345 4.73 1.35 ;
      RECT  4.4 1.35 4.725 1.355 ;
      RECT  4.395 1.355 4.72 1.36 ;
      RECT  4.39 1.36 4.715 1.365 ;
      RECT  4.385 1.365 4.71 1.37 ;
      RECT  4.38 1.37 4.705 1.375 ;
      RECT  4.375 1.375 4.7 1.38 ;
      RECT  4.37 1.38 4.695 1.385 ;
      RECT  4.365 1.385 4.69 1.39 ;
      RECT  4.36 1.39 4.685 1.395 ;
      RECT  4.355 1.395 4.68 1.4 ;
      RECT  4.35 1.4 4.675 1.405 ;
      RECT  4.345 1.405 4.67 1.41 ;
      RECT  4.34 1.41 4.665 1.415 ;
      RECT  4.335 1.415 4.66 1.42 ;
      RECT  4.33 1.42 4.655 1.425 ;
      RECT  4.325 1.425 4.65 1.43 ;
      RECT  4.32 1.43 4.645 1.435 ;
      RECT  4.315 1.435 4.64 1.44 ;
      RECT  4.31 1.44 4.635 1.445 ;
      RECT  4.305 1.445 4.63 1.45 ;
      RECT  4.3 1.45 4.625 1.455 ;
      RECT  4.295 1.455 4.62 1.46 ;
      RECT  4.29 1.46 4.615 1.465 ;
      RECT  4.285 1.465 4.61 1.47 ;
      RECT  4.28 1.47 4.605 1.475 ;
      RECT  4.275 1.475 4.6 1.48 ;
      RECT  4.27 1.48 4.595 1.485 ;
      RECT  4.265 1.485 4.59 1.49 ;
      RECT  4.26 1.49 4.585 1.495 ;
      RECT  4.255 1.495 4.58 1.5 ;
      RECT  4.25 1.5 4.575 1.505 ;
      RECT  4.245 1.505 4.57 1.51 ;
      RECT  4.24 1.51 4.565 1.515 ;
      RECT  4.235 1.515 4.56 1.52 ;
      RECT  4.23 1.52 4.555 1.525 ;
      RECT  4.225 1.525 4.55 1.53 ;
      RECT  4.22 1.53 4.545 1.535 ;
      RECT  4.215 1.535 4.54 1.54 ;
      RECT  4.21 1.54 4.535 1.545 ;
      RECT  4.205 1.545 4.53 1.55 ;
      RECT  4.2 1.55 4.525 1.555 ;
      RECT  4.195 1.555 4.52 1.56 ;
      RECT  4.19 1.56 4.515 1.565 ;
      RECT  1.72 1.565 4.51 1.57 ;
      RECT  1.72 1.57 4.505 1.575 ;
      RECT  1.72 1.575 4.5 1.58 ;
      RECT  1.72 1.58 4.495 1.585 ;
      RECT  1.72 1.585 4.49 1.59 ;
      RECT  1.72 1.59 4.485 1.595 ;
      RECT  1.72 1.595 4.48 1.6 ;
      RECT  1.72 1.6 4.475 1.605 ;
      RECT  1.72 1.605 4.47 1.61 ;
      RECT  1.72 1.61 4.465 1.615 ;
      RECT  1.72 1.615 4.46 1.62 ;
      RECT  1.72 1.62 4.455 1.625 ;
      RECT  1.72 1.625 4.45 1.63 ;
      RECT  1.72 1.63 4.445 1.635 ;
      RECT  1.72 1.635 4.44 1.64 ;
      RECT  1.72 1.64 4.435 1.645 ;
      RECT  1.72 1.645 4.43 1.65 ;
      RECT  1.72 1.65 4.425 1.655 ;
      RECT  1.72 1.655 4.42 1.66 ;
      RECT  1.72 1.66 4.415 1.665 ;
      RECT  1.72 1.665 4.41 1.67 ;
      RECT  1.72 1.67 4.405 1.675 ;
      RECT  1.72 1.675 4.4 1.68 ;
      RECT  1.72 1.68 4.395 1.685 ;
      RECT  1.72 1.685 4.39 1.69 ;
      RECT  1.72 1.69 4.385 1.695 ;
      RECT  1.72 1.695 4.38 1.7 ;
      RECT  1.72 1.7 4.375 1.705 ;
      RECT  1.72 1.705 4.37 1.71 ;
      RECT  1.72 1.71 4.365 1.715 ;
      RECT  1.72 1.715 4.36 1.72 ;
      RECT  1.72 1.72 4.355 1.725 ;
      RECT  1.72 1.725 4.35 1.73 ;
      RECT  1.72 1.73 4.345 1.735 ;
      RECT  1.72 1.735 4.34 1.74 ;
      RECT  1.72 1.74 4.335 1.745 ;
      RECT  1.72 1.745 4.33 1.75 ;
      RECT  1.72 1.75 4.325 1.755 ;
      RECT  1.72 1.755 4.32 1.76 ;
      RECT  1.72 1.76 4.315 1.765 ;
      RECT  1.72 1.765 4.31 1.77 ;
      RECT  1.72 1.77 4.305 1.775 ;
      RECT  1.72 1.775 4.3 1.78 ;
      RECT  1.72 1.78 4.295 1.785 ;
      RECT  1.72 1.785 4.29 1.79 ;
      RECT  1.72 1.79 4.285 1.795 ;
      RECT  12.92 1.29 16.2 1.52 ;
      RECT  8.44 1.565 9.48 1.795 ;
      RECT  12.15 1.565 12.49 1.795 ;
      RECT  12.15 1.795 12.38 3.03 ;
      RECT  12.15 3.03 12.49 3.26 ;
      RECT  11.38 1.75 11.875 1.98 ;
      RECT  11.645 1.98 11.875 3.515 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 3.245 ;
      RECT  6.045 3.245 7.395 3.475 ;
      RECT  7.165 3.475 7.395 3.515 ;
      RECT  7.165 3.515 13.26 3.745 ;
      RECT  9.405 2.35 9.635 3.515 ;
      RECT  13.32 1.75 13.96 1.98 ;
      RECT  13.32 1.98 13.55 2.41 ;
      RECT  12.71 2.41 13.55 2.64 ;
      RECT  13.32 2.64 13.55 3.025 ;
      RECT  13.32 3.025 13.905 3.255 ;
      RECT  13.675 3.255 13.905 4.02 ;
      RECT  10.525 4.02 13.905 4.25 ;
      RECT  10.525 4.25 10.755 4.44 ;
      RECT  9.405 4.44 10.755 4.67 ;
      RECT  9.405 4.67 9.635 5.0 ;
      RECT  7.11 5.0 9.635 5.23 ;
      RECT  14.445 1.75 15.5 1.98 ;
      RECT  14.445 1.98 14.675 2.41 ;
      RECT  13.83 2.41 14.675 2.64 ;
      RECT  14.445 2.64 14.675 3.805 ;
      RECT  14.445 3.805 15.5 4.035 ;
      RECT  4.66 1.75 5.0 2.125 ;
      RECT  3.805 2.125 5.0 2.355 ;
      RECT  3.805 2.355 4.035 3.245 ;
      RECT  3.805 3.245 5.0 3.475 ;
      RECT  1.72 3.805 2.76 4.035 ;
      RECT  6.9 3.975 9.48 4.205 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.925 4.435 8.78 4.665 ;
      RECT  4.925 4.665 5.155 4.925 ;
      RECT  3.19 4.925 5.155 5.155 ;
      RECT  11.38 4.48 16.2 4.71 ;
      RECT  10.47 5.0 12.49 5.23 ;
  END
END MDN_FSDNQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNQ_2
#      Description : D-Flip Flop w/scan, neg-edge triggered, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNQ_2
  CLASS CORE ;
  FOREIGN MDN_FSDNQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.98 2.35 15.26 3.475 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.4 1.565 18.44 1.795 ;
      RECT  17.805 1.795 18.035 3.245 ;
      RECT  17.4 3.245 18.44 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  14.445 4.875 14.675 5.46 ;
      RECT  14.445 5.46 16.915 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  9.965 4.935 10.195 5.46 ;
      RECT  9.965 5.46 11.2 5.74 ;
      RECT  5.485 4.94 5.715 5.46 ;
      RECT  4.48 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 20.33 0.14 ;
      RECT  16.685 0.14 16.915 0.6 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  13.44 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.6 ;
      RECT  9.965 -0.14 11.2 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  4.48 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 4.3 1.12 ;
      RECT  3.245 0.89 4.3 1.005 ;
      RECT  0.18 1.12 3.475 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  18.07 -0.13 18.33 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 5.21 0.6 ;
      RECT  5.99 0.37 7.955 0.6 ;
      RECT  7.725 0.6 7.955 3.315 ;
      RECT  10.455 0.37 14.17 0.6 ;
      RECT  10.455 0.6 10.685 1.005 ;
      RECT  8.23 0.37 8.57 0.6 ;
      RECT  8.23 0.6 8.46 1.005 ;
      RECT  8.23 1.005 10.685 1.235 ;
      RECT  17.185 0.37 18.655 0.6 ;
      RECT  17.185 0.6 17.415 0.83 ;
      RECT  16.07 0.37 16.41 0.6 ;
      RECT  16.18 0.6 16.41 0.83 ;
      RECT  10.915 0.83 17.415 1.06 ;
      RECT  10.915 1.06 11.145 1.565 ;
      RECT  10.525 1.565 11.145 1.795 ;
      RECT  10.525 1.795 10.755 3.03 ;
      RECT  10.525 3.03 11.02 3.26 ;
      RECT  4.745 1.005 7.24 1.01 ;
      RECT  4.74 1.01 7.24 1.015 ;
      RECT  4.735 1.015 7.24 1.02 ;
      RECT  4.73 1.02 7.24 1.025 ;
      RECT  4.725 1.025 7.24 1.03 ;
      RECT  4.72 1.03 7.24 1.035 ;
      RECT  4.715 1.035 7.24 1.04 ;
      RECT  4.71 1.04 7.24 1.045 ;
      RECT  4.705 1.045 7.24 1.05 ;
      RECT  4.7 1.05 7.24 1.055 ;
      RECT  4.695 1.055 7.24 1.06 ;
      RECT  4.69 1.06 7.24 1.065 ;
      RECT  4.685 1.065 7.24 1.07 ;
      RECT  4.68 1.07 7.24 1.075 ;
      RECT  4.675 1.075 7.24 1.08 ;
      RECT  4.67 1.08 7.24 1.085 ;
      RECT  4.665 1.085 7.24 1.09 ;
      RECT  4.66 1.09 7.24 1.095 ;
      RECT  4.655 1.095 7.24 1.1 ;
      RECT  4.65 1.1 7.24 1.105 ;
      RECT  4.645 1.105 7.24 1.11 ;
      RECT  4.64 1.11 7.24 1.115 ;
      RECT  4.635 1.115 7.24 1.12 ;
      RECT  4.63 1.12 7.24 1.125 ;
      RECT  4.625 1.125 7.24 1.13 ;
      RECT  4.62 1.13 7.24 1.135 ;
      RECT  4.615 1.135 7.24 1.14 ;
      RECT  4.61 1.14 7.24 1.145 ;
      RECT  4.605 1.145 7.24 1.15 ;
      RECT  4.6 1.15 7.24 1.155 ;
      RECT  4.595 1.155 7.24 1.16 ;
      RECT  4.59 1.16 7.24 1.165 ;
      RECT  4.585 1.165 7.24 1.17 ;
      RECT  4.58 1.17 7.24 1.175 ;
      RECT  4.575 1.175 7.24 1.18 ;
      RECT  4.57 1.18 7.24 1.185 ;
      RECT  4.565 1.185 7.24 1.19 ;
      RECT  4.56 1.19 7.24 1.195 ;
      RECT  4.555 1.195 7.24 1.2 ;
      RECT  4.55 1.2 7.24 1.205 ;
      RECT  4.545 1.205 7.24 1.21 ;
      RECT  4.54 1.21 7.24 1.215 ;
      RECT  4.535 1.215 7.24 1.22 ;
      RECT  4.53 1.22 7.24 1.225 ;
      RECT  4.525 1.225 7.24 1.23 ;
      RECT  4.52 1.23 7.24 1.235 ;
      RECT  4.515 1.235 4.84 1.24 ;
      RECT  4.51 1.24 4.835 1.245 ;
      RECT  4.505 1.245 4.83 1.25 ;
      RECT  4.5 1.25 4.825 1.255 ;
      RECT  4.495 1.255 4.82 1.26 ;
      RECT  4.49 1.26 4.815 1.265 ;
      RECT  4.485 1.265 4.81 1.27 ;
      RECT  4.48 1.27 4.805 1.275 ;
      RECT  4.475 1.275 4.8 1.28 ;
      RECT  4.47 1.28 4.795 1.285 ;
      RECT  4.465 1.285 4.79 1.29 ;
      RECT  4.46 1.29 4.785 1.295 ;
      RECT  4.455 1.295 4.78 1.3 ;
      RECT  4.45 1.3 4.775 1.305 ;
      RECT  4.445 1.305 4.77 1.31 ;
      RECT  4.44 1.31 4.765 1.315 ;
      RECT  4.435 1.315 4.76 1.32 ;
      RECT  4.43 1.32 4.755 1.325 ;
      RECT  4.425 1.325 4.75 1.33 ;
      RECT  4.42 1.33 4.745 1.335 ;
      RECT  4.415 1.335 4.74 1.34 ;
      RECT  4.41 1.34 4.735 1.345 ;
      RECT  4.405 1.345 4.73 1.35 ;
      RECT  4.4 1.35 4.725 1.355 ;
      RECT  4.395 1.355 4.72 1.36 ;
      RECT  4.39 1.36 4.715 1.365 ;
      RECT  4.385 1.365 4.71 1.37 ;
      RECT  4.38 1.37 4.705 1.375 ;
      RECT  4.375 1.375 4.7 1.38 ;
      RECT  4.37 1.38 4.695 1.385 ;
      RECT  4.365 1.385 4.69 1.39 ;
      RECT  4.36 1.39 4.685 1.395 ;
      RECT  4.355 1.395 4.68 1.4 ;
      RECT  4.35 1.4 4.675 1.405 ;
      RECT  4.345 1.405 4.67 1.41 ;
      RECT  4.34 1.41 4.665 1.415 ;
      RECT  4.335 1.415 4.66 1.42 ;
      RECT  4.33 1.42 4.655 1.425 ;
      RECT  4.325 1.425 4.65 1.43 ;
      RECT  4.32 1.43 4.645 1.435 ;
      RECT  4.315 1.435 4.64 1.44 ;
      RECT  4.31 1.44 4.635 1.445 ;
      RECT  4.305 1.445 4.63 1.45 ;
      RECT  4.3 1.45 4.625 1.455 ;
      RECT  4.295 1.455 4.62 1.46 ;
      RECT  4.29 1.46 4.615 1.465 ;
      RECT  4.285 1.465 4.61 1.47 ;
      RECT  4.28 1.47 4.605 1.475 ;
      RECT  4.275 1.475 4.6 1.48 ;
      RECT  4.27 1.48 4.595 1.485 ;
      RECT  4.265 1.485 4.59 1.49 ;
      RECT  4.26 1.49 4.585 1.495 ;
      RECT  4.255 1.495 4.58 1.5 ;
      RECT  4.25 1.5 4.575 1.505 ;
      RECT  4.245 1.505 4.57 1.51 ;
      RECT  4.24 1.51 4.565 1.515 ;
      RECT  4.235 1.515 4.56 1.52 ;
      RECT  4.23 1.52 4.555 1.525 ;
      RECT  4.225 1.525 4.55 1.53 ;
      RECT  4.22 1.53 4.545 1.535 ;
      RECT  4.215 1.535 4.54 1.54 ;
      RECT  4.21 1.54 4.535 1.545 ;
      RECT  4.205 1.545 4.53 1.55 ;
      RECT  4.2 1.55 4.525 1.555 ;
      RECT  4.195 1.555 4.52 1.56 ;
      RECT  4.19 1.56 4.515 1.565 ;
      RECT  1.72 1.565 4.51 1.57 ;
      RECT  1.72 1.57 4.505 1.575 ;
      RECT  1.72 1.575 4.5 1.58 ;
      RECT  1.72 1.58 4.495 1.585 ;
      RECT  1.72 1.585 4.49 1.59 ;
      RECT  1.72 1.59 4.485 1.595 ;
      RECT  1.72 1.595 4.48 1.6 ;
      RECT  1.72 1.6 4.475 1.605 ;
      RECT  1.72 1.605 4.47 1.61 ;
      RECT  1.72 1.61 4.465 1.615 ;
      RECT  1.72 1.615 4.46 1.62 ;
      RECT  1.72 1.62 4.455 1.625 ;
      RECT  1.72 1.625 4.45 1.63 ;
      RECT  1.72 1.63 4.445 1.635 ;
      RECT  1.72 1.635 4.44 1.64 ;
      RECT  1.72 1.64 4.435 1.645 ;
      RECT  1.72 1.645 4.43 1.65 ;
      RECT  1.72 1.65 4.425 1.655 ;
      RECT  1.72 1.655 4.42 1.66 ;
      RECT  1.72 1.66 4.415 1.665 ;
      RECT  1.72 1.665 4.41 1.67 ;
      RECT  1.72 1.67 4.405 1.675 ;
      RECT  1.72 1.675 4.4 1.68 ;
      RECT  1.72 1.68 4.395 1.685 ;
      RECT  1.72 1.685 4.39 1.69 ;
      RECT  1.72 1.69 4.385 1.695 ;
      RECT  1.72 1.695 4.38 1.7 ;
      RECT  1.72 1.7 4.375 1.705 ;
      RECT  1.72 1.705 4.37 1.71 ;
      RECT  1.72 1.71 4.365 1.715 ;
      RECT  1.72 1.715 4.36 1.72 ;
      RECT  1.72 1.72 4.355 1.725 ;
      RECT  1.72 1.725 4.35 1.73 ;
      RECT  1.72 1.73 4.345 1.735 ;
      RECT  1.72 1.735 4.34 1.74 ;
      RECT  1.72 1.74 4.335 1.745 ;
      RECT  1.72 1.745 4.33 1.75 ;
      RECT  1.72 1.75 4.325 1.755 ;
      RECT  1.72 1.755 4.32 1.76 ;
      RECT  1.72 1.76 4.315 1.765 ;
      RECT  1.72 1.765 4.31 1.77 ;
      RECT  1.72 1.77 4.305 1.775 ;
      RECT  1.72 1.775 4.3 1.78 ;
      RECT  1.72 1.78 4.295 1.785 ;
      RECT  1.72 1.785 4.29 1.79 ;
      RECT  1.72 1.79 4.285 1.795 ;
      RECT  12.92 1.29 16.2 1.52 ;
      RECT  8.44 1.565 9.48 1.795 ;
      RECT  11.38 1.565 11.875 1.795 ;
      RECT  11.645 1.795 11.875 3.49 ;
      RECT  9.405 2.35 9.635 3.245 ;
      RECT  8.285 3.245 9.635 3.475 ;
      RECT  9.405 3.475 9.635 3.49 ;
      RECT  8.285 3.475 8.515 3.545 ;
      RECT  9.405 3.49 13.26 3.71 ;
      RECT  12.92 3.48 13.26 3.49 ;
      RECT  6.255 1.51 6.485 3.545 ;
      RECT  6.25 3.545 8.515 3.775 ;
      RECT  9.405 3.71 13.11 3.72 ;
      RECT  12.15 1.565 12.49 1.795 ;
      RECT  12.15 1.795 12.38 3.03 ;
      RECT  12.15 3.03 12.49 3.26 ;
      RECT  13.325 1.75 13.96 1.98 ;
      RECT  13.325 1.98 13.555 2.405 ;
      RECT  12.71 2.405 13.555 2.635 ;
      RECT  13.325 2.635 13.555 3.025 ;
      RECT  13.325 3.025 14.12 3.255 ;
      RECT  13.89 3.255 14.12 3.95 ;
      RECT  10.525 3.95 14.12 4.18 ;
      RECT  10.525 4.18 10.755 4.475 ;
      RECT  9.405 4.475 10.755 4.705 ;
      RECT  9.405 4.705 9.635 5.0 ;
      RECT  7.11 5.0 9.635 5.23 ;
      RECT  14.445 1.75 15.5 1.98 ;
      RECT  14.445 1.98 14.675 2.405 ;
      RECT  13.83 2.405 14.675 2.635 ;
      RECT  14.445 2.635 14.675 3.805 ;
      RECT  14.445 3.805 15.5 4.035 ;
      RECT  4.715 1.695 4.945 2.125 ;
      RECT  3.805 2.125 5.715 2.355 ;
      RECT  3.805 2.355 4.035 2.69 ;
      RECT  5.485 2.355 5.715 3.805 ;
      RECT  4.66 3.805 5.715 4.035 ;
      RECT  1.72 3.805 2.76 4.035 ;
      RECT  6.9 4.015 9.48 4.245 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  11.38 4.415 16.2 4.645 ;
      RECT  4.925 4.48 8.78 4.71 ;
      RECT  4.925 4.71 5.155 4.985 ;
      RECT  3.19 4.985 5.155 5.215 ;
      RECT  10.47 5.0 12.49 5.23 ;
  END
END MDN_FSDNQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNQ_4
#      Description : D-Flip Flop w/scan, neg-edge triggered, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNQ_4
  CLASS CORE ;
  FOREIGN MDN_FSDNQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.98 2.35 15.26 3.475 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.4 1.565 20.68 1.795 ;
      RECT  18.925 1.795 19.155 3.245 ;
      RECT  17.4 3.245 20.68 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  14.445 4.94 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  9.965 4.975 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  5.485 4.94 5.715 5.46 ;
      RECT  4.48 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.595 ;
      RECT  13.44 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.595 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.52 ;
      RECT  4.48 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 4.3 1.12 ;
      RECT  3.805 0.89 4.3 1.005 ;
      RECT  0.18 1.12 4.035 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  20.31 -0.13 20.57 0.13 ;
      RECT  20.87 -0.13 21.13 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 5.21 0.6 ;
      RECT  5.99 0.37 7.955 0.6 ;
      RECT  7.725 0.6 7.955 3.315 ;
      RECT  10.525 0.37 14.17 0.6 ;
      RECT  10.525 0.6 10.755 0.785 ;
      RECT  8.23 0.37 8.57 0.6 ;
      RECT  8.34 0.6 8.57 0.785 ;
      RECT  8.34 0.785 10.755 1.015 ;
      RECT  19.43 0.37 20.89 0.6 ;
      RECT  19.43 0.6 19.66 1.005 ;
      RECT  17.19 0.37 18.65 0.6 ;
      RECT  17.19 0.6 17.42 0.83 ;
      RECT  18.42 0.6 18.65 1.005 ;
      RECT  16.07 0.37 16.41 0.6 ;
      RECT  16.18 0.6 16.41 0.83 ;
      RECT  11.085 0.83 17.42 1.06 ;
      RECT  18.42 1.005 19.66 1.235 ;
      RECT  11.085 1.06 11.315 1.295 ;
      RECT  10.525 1.295 11.315 1.525 ;
      RECT  10.525 1.525 10.755 3.03 ;
      RECT  10.525 3.03 11.02 3.26 ;
      RECT  4.745 1.005 7.24 1.01 ;
      RECT  4.74 1.01 7.24 1.015 ;
      RECT  4.735 1.015 7.24 1.02 ;
      RECT  4.73 1.02 7.24 1.025 ;
      RECT  4.725 1.025 7.24 1.03 ;
      RECT  4.72 1.03 7.24 1.035 ;
      RECT  4.715 1.035 7.24 1.04 ;
      RECT  4.71 1.04 7.24 1.045 ;
      RECT  4.705 1.045 7.24 1.05 ;
      RECT  4.7 1.05 7.24 1.055 ;
      RECT  4.695 1.055 7.24 1.06 ;
      RECT  4.69 1.06 7.24 1.065 ;
      RECT  4.685 1.065 7.24 1.07 ;
      RECT  4.68 1.07 7.24 1.075 ;
      RECT  4.675 1.075 7.24 1.08 ;
      RECT  4.67 1.08 7.24 1.085 ;
      RECT  4.665 1.085 7.24 1.09 ;
      RECT  4.66 1.09 7.24 1.095 ;
      RECT  4.655 1.095 7.24 1.1 ;
      RECT  4.65 1.1 7.24 1.105 ;
      RECT  4.645 1.105 7.24 1.11 ;
      RECT  4.64 1.11 7.24 1.115 ;
      RECT  4.635 1.115 7.24 1.12 ;
      RECT  4.63 1.12 7.24 1.125 ;
      RECT  4.625 1.125 7.24 1.13 ;
      RECT  4.62 1.13 7.24 1.135 ;
      RECT  4.615 1.135 7.24 1.14 ;
      RECT  4.61 1.14 7.24 1.145 ;
      RECT  4.605 1.145 7.24 1.15 ;
      RECT  4.6 1.15 7.24 1.155 ;
      RECT  4.595 1.155 7.24 1.16 ;
      RECT  4.59 1.16 7.24 1.165 ;
      RECT  4.585 1.165 7.24 1.17 ;
      RECT  4.58 1.17 7.24 1.175 ;
      RECT  4.575 1.175 7.24 1.18 ;
      RECT  4.57 1.18 7.24 1.185 ;
      RECT  4.565 1.185 7.24 1.19 ;
      RECT  4.56 1.19 7.24 1.195 ;
      RECT  4.555 1.195 7.24 1.2 ;
      RECT  4.55 1.2 7.24 1.205 ;
      RECT  4.545 1.205 7.24 1.21 ;
      RECT  4.54 1.21 7.24 1.215 ;
      RECT  4.535 1.215 7.24 1.22 ;
      RECT  4.53 1.22 7.24 1.225 ;
      RECT  4.525 1.225 7.24 1.23 ;
      RECT  4.52 1.23 7.24 1.235 ;
      RECT  4.515 1.235 4.84 1.24 ;
      RECT  4.51 1.24 4.835 1.245 ;
      RECT  4.505 1.245 4.83 1.25 ;
      RECT  4.5 1.25 4.825 1.255 ;
      RECT  4.495 1.255 4.82 1.26 ;
      RECT  4.49 1.26 4.815 1.265 ;
      RECT  4.485 1.265 4.81 1.27 ;
      RECT  4.48 1.27 4.805 1.275 ;
      RECT  4.475 1.275 4.8 1.28 ;
      RECT  4.47 1.28 4.795 1.285 ;
      RECT  4.465 1.285 4.79 1.29 ;
      RECT  4.46 1.29 4.785 1.295 ;
      RECT  4.455 1.295 4.78 1.3 ;
      RECT  4.45 1.3 4.775 1.305 ;
      RECT  4.445 1.305 4.77 1.31 ;
      RECT  4.44 1.31 4.765 1.315 ;
      RECT  4.435 1.315 4.76 1.32 ;
      RECT  4.43 1.32 4.755 1.325 ;
      RECT  4.425 1.325 4.75 1.33 ;
      RECT  4.42 1.33 4.745 1.335 ;
      RECT  4.415 1.335 4.74 1.34 ;
      RECT  4.41 1.34 4.735 1.345 ;
      RECT  4.405 1.345 4.73 1.35 ;
      RECT  4.4 1.35 4.725 1.355 ;
      RECT  4.395 1.355 4.72 1.36 ;
      RECT  4.39 1.36 4.715 1.365 ;
      RECT  4.385 1.365 4.71 1.37 ;
      RECT  4.38 1.37 4.705 1.375 ;
      RECT  4.375 1.375 4.7 1.38 ;
      RECT  4.37 1.38 4.695 1.385 ;
      RECT  4.365 1.385 4.69 1.39 ;
      RECT  4.36 1.39 4.685 1.395 ;
      RECT  4.355 1.395 4.68 1.4 ;
      RECT  4.35 1.4 4.675 1.405 ;
      RECT  4.345 1.405 4.67 1.41 ;
      RECT  4.34 1.41 4.665 1.415 ;
      RECT  4.335 1.415 4.66 1.42 ;
      RECT  4.33 1.42 4.655 1.425 ;
      RECT  4.325 1.425 4.65 1.43 ;
      RECT  4.32 1.43 4.645 1.435 ;
      RECT  4.315 1.435 4.64 1.44 ;
      RECT  4.31 1.44 4.635 1.445 ;
      RECT  4.305 1.445 4.63 1.45 ;
      RECT  4.3 1.45 4.625 1.455 ;
      RECT  4.295 1.455 4.62 1.46 ;
      RECT  4.29 1.46 4.615 1.465 ;
      RECT  4.285 1.465 4.61 1.47 ;
      RECT  4.28 1.47 4.605 1.475 ;
      RECT  4.275 1.475 4.6 1.48 ;
      RECT  4.27 1.48 4.595 1.485 ;
      RECT  4.265 1.485 4.59 1.49 ;
      RECT  4.26 1.49 4.585 1.495 ;
      RECT  4.255 1.495 4.58 1.5 ;
      RECT  4.25 1.5 4.575 1.505 ;
      RECT  4.245 1.505 4.57 1.51 ;
      RECT  4.24 1.51 4.565 1.515 ;
      RECT  4.235 1.515 4.56 1.52 ;
      RECT  4.23 1.52 4.555 1.525 ;
      RECT  4.225 1.525 4.55 1.53 ;
      RECT  4.22 1.53 4.545 1.535 ;
      RECT  4.215 1.535 4.54 1.54 ;
      RECT  4.21 1.54 4.535 1.545 ;
      RECT  4.205 1.545 4.53 1.55 ;
      RECT  4.2 1.55 4.525 1.555 ;
      RECT  4.195 1.555 4.52 1.56 ;
      RECT  4.19 1.56 4.515 1.565 ;
      RECT  1.72 1.565 4.51 1.57 ;
      RECT  1.72 1.57 4.505 1.575 ;
      RECT  1.72 1.575 4.5 1.58 ;
      RECT  1.72 1.58 4.495 1.585 ;
      RECT  1.72 1.585 4.49 1.59 ;
      RECT  1.72 1.59 4.485 1.595 ;
      RECT  1.72 1.595 4.48 1.6 ;
      RECT  1.72 1.6 4.475 1.605 ;
      RECT  1.72 1.605 4.47 1.61 ;
      RECT  1.72 1.61 4.465 1.615 ;
      RECT  1.72 1.615 4.46 1.62 ;
      RECT  1.72 1.62 4.455 1.625 ;
      RECT  1.72 1.625 4.45 1.63 ;
      RECT  1.72 1.63 4.445 1.635 ;
      RECT  1.72 1.635 4.44 1.64 ;
      RECT  1.72 1.64 4.435 1.645 ;
      RECT  1.72 1.645 4.43 1.65 ;
      RECT  1.72 1.65 4.425 1.655 ;
      RECT  1.72 1.655 4.42 1.66 ;
      RECT  1.72 1.66 4.415 1.665 ;
      RECT  1.72 1.665 4.41 1.67 ;
      RECT  1.72 1.67 4.405 1.675 ;
      RECT  1.72 1.675 4.4 1.68 ;
      RECT  1.72 1.68 4.395 1.685 ;
      RECT  1.72 1.685 4.39 1.69 ;
      RECT  1.72 1.69 4.385 1.695 ;
      RECT  1.72 1.695 4.38 1.7 ;
      RECT  1.72 1.7 4.375 1.705 ;
      RECT  1.72 1.705 4.37 1.71 ;
      RECT  1.72 1.71 4.365 1.715 ;
      RECT  1.72 1.715 4.36 1.72 ;
      RECT  1.72 1.72 4.355 1.725 ;
      RECT  1.72 1.725 4.35 1.73 ;
      RECT  1.72 1.73 4.345 1.735 ;
      RECT  1.72 1.735 4.34 1.74 ;
      RECT  1.72 1.74 4.335 1.745 ;
      RECT  1.72 1.745 4.33 1.75 ;
      RECT  1.72 1.75 4.325 1.755 ;
      RECT  1.72 1.755 4.32 1.76 ;
      RECT  1.72 1.76 4.315 1.765 ;
      RECT  1.72 1.765 4.31 1.77 ;
      RECT  1.72 1.77 4.305 1.775 ;
      RECT  1.72 1.775 4.3 1.78 ;
      RECT  1.72 1.78 4.295 1.785 ;
      RECT  1.72 1.785 4.29 1.79 ;
      RECT  1.72 1.79 4.285 1.795 ;
      RECT  12.92 1.29 16.2 1.52 ;
      RECT  8.44 1.565 9.48 1.795 ;
      RECT  4.66 1.75 5.155 1.98 ;
      RECT  4.925 1.98 5.155 2.685 ;
      RECT  3.805 2.345 4.035 2.685 ;
      RECT  3.805 2.685 5.155 2.915 ;
      RECT  4.925 2.915 5.155 3.805 ;
      RECT  4.66 3.805 5.155 4.035 ;
      RECT  11.38 1.75 11.875 1.98 ;
      RECT  11.645 1.98 11.875 3.545 ;
      RECT  6.255 1.51 6.485 3.545 ;
      RECT  6.255 3.545 13.26 3.775 ;
      RECT  9.405 2.35 9.635 3.545 ;
      RECT  13.325 1.75 13.96 1.98 ;
      RECT  13.325 1.98 13.555 2.405 ;
      RECT  12.71 2.405 13.555 2.635 ;
      RECT  13.325 2.635 13.555 3.025 ;
      RECT  13.325 3.025 13.905 3.255 ;
      RECT  13.675 3.255 13.905 4.02 ;
      RECT  10.525 4.02 13.905 4.25 ;
      RECT  10.525 4.25 10.755 4.515 ;
      RECT  9.405 4.515 10.755 4.745 ;
      RECT  9.405 4.745 9.635 5.0 ;
      RECT  7.11 5.0 9.635 5.23 ;
      RECT  14.445 1.75 15.5 1.98 ;
      RECT  14.445 1.98 14.675 2.405 ;
      RECT  13.83 2.405 14.675 2.635 ;
      RECT  14.445 2.635 14.675 3.805 ;
      RECT  14.445 3.805 15.5 4.035 ;
      RECT  12.205 1.51 12.435 3.315 ;
      RECT  1.72 3.805 2.76 4.035 ;
      RECT  6.9 4.015 9.48 4.245 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.925 4.475 8.78 4.705 ;
      RECT  4.925 4.705 5.155 4.925 ;
      RECT  3.19 4.925 5.155 5.155 ;
      RECT  11.38 4.48 16.2 4.71 ;
      RECT  10.47 5.0 12.49 5.23 ;
  END
END MDN_FSDNQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNRB_4
#      Description : D-Flip Flop w/scan, neg-edge triggered, lo-async-clear
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNRB_4
  CLASS CORE ;
  FOREIGN MDN_FSDNRB_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 29.12 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 1.565 2.94 2.69 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.64 1.565 22.92 1.795 ;
      RECT  22.285 1.795 22.515 3.245 ;
      RECT  19.64 3.245 22.92 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  24.82 1.565 28.94 1.795 ;
      RECT  26.765 1.795 26.995 3.245 ;
      RECT  24.82 3.245 28.94 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END QN
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.98 2.125 16.38 2.355 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  27.885 4.9 28.115 5.46 ;
      RECT  27.885 5.46 29.29 5.74 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.645 5.46 26.32 5.74 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.08 5.74 ;
      RECT  21.165 4.905 21.395 5.46 ;
      RECT  20.72 5.46 21.395 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  14.445 5.08 14.675 5.46 ;
      RECT  13.27 5.46 15.12 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 11.2 5.74 ;
      RECT  5.43 5.135 5.77 5.46 ;
      RECT  5.04 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 29.12 5.74 ;
      LAYER VIA12 ;
      RECT  28.15 5.47 28.41 5.73 ;
      RECT  28.71 5.47 28.97 5.73 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 -0.14 29.29 0.14 ;
      RECT  25.645 0.14 25.875 0.7 ;
      RECT  27.885 0.14 28.115 0.7 ;
      RECT  21.16 -0.14 23.635 0.14 ;
      RECT  21.16 0.14 21.4 0.7 ;
      RECT  23.405 0.14 23.635 0.73 ;
      RECT  18.48 -0.14 19.16 0.14 ;
      RECT  18.92 0.14 19.16 0.7 ;
      RECT  15.12 -0.14 16.24 0.14 ;
      RECT  15.565 0.14 15.795 0.89 ;
      RECT  15.16 0.89 16.2 1.12 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.52 ;
      RECT  3.805 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.52 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 29.12 0.14 ;
      LAYER VIA12 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  27.03 -0.13 27.29 0.13 ;
      RECT  27.59 -0.13 27.85 0.13 ;
      RECT  28.15 -0.13 28.41 0.13 ;
      RECT  28.71 -0.13 28.97 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  22.55 -0.13 22.81 0.13 ;
      RECT  23.11 -0.13 23.37 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  10.515 0.37 13.05 0.6 ;
      RECT  10.515 0.6 10.745 0.75 ;
      RECT  5.98 0.37 9.635 0.6 ;
      RECT  5.98 0.6 6.21 0.75 ;
      RECT  9.405 0.6 9.635 0.75 ;
      RECT  4.66 0.75 6.21 0.98 ;
      RECT  9.405 0.75 10.745 0.98 ;
      RECT  4.66 0.98 5.0 1.12 ;
      RECT  23.91 0.37 24.25 0.6 ;
      RECT  23.91 0.6 24.14 1.005 ;
      RECT  21.67 0.37 23.13 0.6 ;
      RECT  22.845 0.6 23.075 1.005 ;
      RECT  22.845 1.005 24.14 1.235 ;
      RECT  26.15 0.37 27.61 0.6 ;
      RECT  6.44 0.83 8.78 1.06 ;
      RECT  8.44 1.06 8.78 1.12 ;
      RECT  6.44 1.06 6.67 1.215 ;
      RECT  5.225 1.215 6.67 1.445 ;
      RECT  5.225 1.445 5.455 1.565 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  3.245 1.565 5.455 1.795 ;
      RECT  10.975 0.83 13.96 1.06 ;
      RECT  13.62 1.06 13.96 1.12 ;
      RECT  10.975 1.06 11.205 1.29 ;
      RECT  8.945 1.29 11.205 1.295 ;
      RECT  8.94 1.295 11.205 1.3 ;
      RECT  8.935 1.3 11.205 1.305 ;
      RECT  8.93 1.305 11.205 1.31 ;
      RECT  8.925 1.31 11.205 1.315 ;
      RECT  8.92 1.315 11.205 1.32 ;
      RECT  8.915 1.32 11.205 1.325 ;
      RECT  8.91 1.325 11.205 1.33 ;
      RECT  8.905 1.33 11.205 1.335 ;
      RECT  8.9 1.335 11.205 1.34 ;
      RECT  8.895 1.34 11.205 1.345 ;
      RECT  8.89 1.345 11.205 1.35 ;
      RECT  6.9 1.29 8.215 1.295 ;
      RECT  6.9 1.295 8.22 1.3 ;
      RECT  6.9 1.3 8.225 1.305 ;
      RECT  6.9 1.305 8.23 1.31 ;
      RECT  6.9 1.31 8.235 1.315 ;
      RECT  6.9 1.315 8.24 1.32 ;
      RECT  6.9 1.32 8.245 1.325 ;
      RECT  6.9 1.325 8.25 1.33 ;
      RECT  6.9 1.33 8.255 1.335 ;
      RECT  6.9 1.335 8.26 1.34 ;
      RECT  6.9 1.34 8.265 1.345 ;
      RECT  6.9 1.345 8.27 1.35 ;
      RECT  6.9 1.35 11.205 1.52 ;
      RECT  8.11 1.52 9.04 1.525 ;
      RECT  8.115 1.525 9.035 1.53 ;
      RECT  8.12 1.53 9.03 1.535 ;
      RECT  8.125 1.535 9.025 1.54 ;
      RECT  8.13 1.54 9.02 1.545 ;
      RECT  8.135 1.545 9.015 1.55 ;
      RECT  8.14 1.55 9.01 1.555 ;
      RECT  8.145 1.555 9.005 1.56 ;
      RECT  8.15 1.56 9.0 1.565 ;
      RECT  8.155 1.565 8.995 1.57 ;
      RECT  8.16 1.57 8.99 1.575 ;
      RECT  8.165 1.575 8.985 1.58 ;
      RECT  16.685 1.005 18.44 1.235 ;
      RECT  16.685 1.235 16.915 1.35 ;
      RECT  11.435 1.29 13.46 1.295 ;
      RECT  11.435 1.295 13.465 1.3 ;
      RECT  11.435 1.3 13.47 1.305 ;
      RECT  11.435 1.305 13.475 1.31 ;
      RECT  11.435 1.31 13.48 1.315 ;
      RECT  11.435 1.315 13.485 1.32 ;
      RECT  11.435 1.32 13.49 1.325 ;
      RECT  11.435 1.325 13.495 1.33 ;
      RECT  11.435 1.33 13.5 1.335 ;
      RECT  11.435 1.335 13.505 1.34 ;
      RECT  11.435 1.34 13.51 1.345 ;
      RECT  11.435 1.345 13.515 1.35 ;
      RECT  11.435 1.35 16.915 1.52 ;
      RECT  13.355 1.52 16.915 1.525 ;
      RECT  11.435 1.52 11.665 1.67 ;
      RECT  13.36 1.525 16.915 1.53 ;
      RECT  13.365 1.53 16.915 1.535 ;
      RECT  13.37 1.535 16.915 1.54 ;
      RECT  13.375 1.54 16.915 1.545 ;
      RECT  13.38 1.545 16.915 1.55 ;
      RECT  13.385 1.55 16.915 1.555 ;
      RECT  13.39 1.555 16.915 1.56 ;
      RECT  13.395 1.56 16.915 1.565 ;
      RECT  13.4 1.565 16.915 1.57 ;
      RECT  13.405 1.57 16.915 1.575 ;
      RECT  13.41 1.575 16.915 1.58 ;
      RECT  17.4 1.565 18.595 1.795 ;
      RECT  18.365 1.795 18.595 2.405 ;
      RECT  18.365 2.405 21.89 2.635 ;
      RECT  18.365 2.635 18.595 3.245 ;
      RECT  15.86 3.245 18.595 3.475 ;
      RECT  23.965 1.565 24.46 1.795 ;
      RECT  23.965 1.795 24.195 2.405 ;
      RECT  23.965 2.405 26.395 2.635 ;
      RECT  23.965 2.635 24.195 3.245 ;
      RECT  23.965 3.245 24.46 3.475 ;
      RECT  7.67 1.75 8.01 1.81 ;
      RECT  7.67 1.81 8.86 2.04 ;
      RECT  8.63 2.04 8.86 2.66 ;
      RECT  8.63 2.66 9.15 2.895 ;
      RECT  7.725 2.895 9.15 2.94 ;
      RECT  7.725 2.94 8.86 3.125 ;
      RECT  7.725 3.125 7.955 3.53 ;
      RECT  6.2 1.675 6.565 1.905 ;
      RECT  6.335 1.905 6.565 2.415 ;
      RECT  6.335 2.415 8.345 2.645 ;
      RECT  6.335 2.645 6.565 3.09 ;
      RECT  6.2 3.09 6.565 3.32 ;
      RECT  9.14 1.75 10.195 1.98 ;
      RECT  9.965 1.98 10.195 3.755 ;
      RECT  8.285 3.755 10.195 3.985 ;
      RECT  8.285 3.985 8.515 4.02 ;
      RECT  7.725 4.02 8.515 4.25 ;
      RECT  7.725 4.25 7.955 4.995 ;
      RECT  4.925 4.675 6.275 4.905 ;
      RECT  6.045 4.905 6.275 4.995 ;
      RECT  4.925 4.905 5.155 5.0 ;
      RECT  6.045 4.995 7.955 5.225 ;
      RECT  3.75 5.0 5.155 5.23 ;
      RECT  12.15 1.75 12.49 1.98 ;
      RECT  12.205 1.98 12.435 3.315 ;
      RECT  12.765 1.75 13.26 1.98 ;
      RECT  12.765 1.98 12.995 2.41 ;
      RECT  12.765 2.41 14.17 2.635 ;
      RECT  13.83 2.405 14.17 2.41 ;
      RECT  12.765 2.635 14.165 2.64 ;
      RECT  12.765 2.64 12.995 3.32 ;
      RECT  12.76 3.32 12.995 3.325 ;
      RECT  12.755 3.325 12.995 3.33 ;
      RECT  12.75 3.33 12.995 3.335 ;
      RECT  12.745 3.335 12.995 3.34 ;
      RECT  12.74 3.34 12.995 3.345 ;
      RECT  12.735 3.345 12.995 3.35 ;
      RECT  12.73 3.35 12.995 3.355 ;
      RECT  12.725 3.355 12.995 3.36 ;
      RECT  12.72 3.36 12.995 3.365 ;
      RECT  12.715 3.365 12.995 3.37 ;
      RECT  12.71 3.37 12.995 3.375 ;
      RECT  12.705 3.375 12.995 3.38 ;
      RECT  12.7 3.38 12.995 3.385 ;
      RECT  12.695 3.385 12.995 3.39 ;
      RECT  12.69 3.39 12.995 3.395 ;
      RECT  12.685 3.395 12.995 3.4 ;
      RECT  12.68 3.4 12.995 3.405 ;
      RECT  12.675 3.405 12.995 3.41 ;
      RECT  12.67 3.41 12.995 3.415 ;
      RECT  12.665 3.415 12.99 3.42 ;
      RECT  12.66 3.42 12.985 3.425 ;
      RECT  12.655 3.425 12.98 3.43 ;
      RECT  12.65 3.43 12.975 3.435 ;
      RECT  12.645 3.435 12.97 3.44 ;
      RECT  12.64 3.44 12.965 3.445 ;
      RECT  12.635 3.445 12.96 3.45 ;
      RECT  12.63 3.45 12.955 3.455 ;
      RECT  12.625 3.455 12.95 3.46 ;
      RECT  12.62 3.46 12.945 3.465 ;
      RECT  12.615 3.465 12.94 3.47 ;
      RECT  12.61 3.47 12.935 3.475 ;
      RECT  12.605 3.475 12.93 3.48 ;
      RECT  12.6 3.48 12.925 3.485 ;
      RECT  12.595 3.485 12.92 3.49 ;
      RECT  12.59 3.49 12.915 3.495 ;
      RECT  12.585 3.495 12.91 3.5 ;
      RECT  12.58 3.5 12.905 3.505 ;
      RECT  12.575 3.505 12.9 3.51 ;
      RECT  12.57 3.51 12.895 3.515 ;
      RECT  12.565 3.515 12.89 3.52 ;
      RECT  12.56 3.52 12.885 3.525 ;
      RECT  12.555 3.525 12.88 3.53 ;
      RECT  12.55 3.53 12.875 3.535 ;
      RECT  12.545 3.535 12.87 3.54 ;
      RECT  12.54 3.54 12.865 3.545 ;
      RECT  12.535 3.545 12.86 3.55 ;
      RECT  10.68 1.75 11.02 1.9 ;
      RECT  10.68 1.9 11.315 2.13 ;
      RECT  11.085 2.13 11.315 3.55 ;
      RECT  10.68 3.55 12.855 3.555 ;
      RECT  10.68 3.555 12.85 3.56 ;
      RECT  10.68 3.56 12.845 3.565 ;
      RECT  10.68 3.565 12.84 3.57 ;
      RECT  10.68 3.57 12.835 3.575 ;
      RECT  10.68 3.575 12.83 3.58 ;
      RECT  10.68 3.58 12.825 3.585 ;
      RECT  10.68 3.585 12.82 3.59 ;
      RECT  10.68 3.59 12.815 3.595 ;
      RECT  10.68 3.595 12.81 3.6 ;
      RECT  10.68 3.6 12.805 3.605 ;
      RECT  10.68 3.605 12.8 3.61 ;
      RECT  10.68 3.61 12.795 3.615 ;
      RECT  10.68 3.615 12.79 3.62 ;
      RECT  10.68 3.62 12.785 3.625 ;
      RECT  10.68 3.625 12.78 3.63 ;
      RECT  10.68 3.63 12.775 3.635 ;
      RECT  10.68 3.635 12.77 3.64 ;
      RECT  10.68 3.64 12.765 3.645 ;
      RECT  10.68 3.645 12.76 3.65 ;
      RECT  10.68 3.65 12.755 3.655 ;
      RECT  10.68 3.655 12.75 3.66 ;
      RECT  10.68 3.66 12.745 3.665 ;
      RECT  10.68 3.665 12.74 3.67 ;
      RECT  10.68 3.67 12.735 3.675 ;
      RECT  10.68 3.675 12.73 3.68 ;
      RECT  10.68 3.68 12.725 3.685 ;
      RECT  10.68 3.685 12.72 3.69 ;
      RECT  10.68 3.69 12.715 3.695 ;
      RECT  10.68 3.695 12.71 3.7 ;
      RECT  10.68 3.7 12.705 3.705 ;
      RECT  10.68 3.705 12.7 3.71 ;
      RECT  10.68 3.71 12.695 3.715 ;
      RECT  10.68 3.715 12.69 3.72 ;
      RECT  10.68 3.72 12.685 3.725 ;
      RECT  10.68 3.725 12.68 3.73 ;
      RECT  10.68 3.73 12.675 3.735 ;
      RECT  10.68 3.735 12.67 3.74 ;
      RECT  10.68 3.74 12.665 3.745 ;
      RECT  10.68 3.745 12.66 3.75 ;
      RECT  10.68 3.75 12.655 3.755 ;
      RECT  10.68 3.755 12.65 3.76 ;
      RECT  10.68 3.76 12.645 3.765 ;
      RECT  10.68 3.765 12.64 3.77 ;
      RECT  10.68 3.77 12.635 3.775 ;
      RECT  10.68 3.775 12.63 3.78 ;
      RECT  27.27 2.405 28.73 2.635 ;
      RECT  5.485 2.445 6.105 2.675 ;
      RECT  5.485 2.675 5.715 3.245 ;
      RECT  4.66 3.245 5.715 3.475 ;
      RECT  10.45 2.36 10.83 2.94 ;
      RECT  9.405 2.345 9.635 3.22 ;
      RECT  9.17 3.22 9.635 3.5 ;
      RECT  1.72 3.145 2.76 3.375 ;
      RECT  3.245 3.245 4.3 3.475 ;
      RECT  3.245 3.475 3.475 3.605 ;
      RECT  2.125 3.605 3.475 3.835 ;
      RECT  2.125 3.835 2.355 4.365 ;
      RECT  0.18 4.365 2.355 4.595 ;
      RECT  7.115 3.22 7.495 3.5 ;
      RECT  7.115 3.5 7.345 3.755 ;
      RECT  3.805 3.755 7.345 3.985 ;
      RECT  3.805 3.985 4.035 4.065 ;
      RECT  2.685 4.065 4.035 4.295 ;
      RECT  2.685 4.295 2.915 5.0 ;
      RECT  1.51 5.0 2.915 5.23 ;
      RECT  13.055 3.685 15.5 3.69 ;
      RECT  13.05 3.69 15.5 3.695 ;
      RECT  13.045 3.695 15.5 3.7 ;
      RECT  13.04 3.7 15.5 3.705 ;
      RECT  13.035 3.705 15.5 3.71 ;
      RECT  13.03 3.71 15.5 3.715 ;
      RECT  13.025 3.715 15.5 3.72 ;
      RECT  13.02 3.72 15.5 3.725 ;
      RECT  13.015 3.725 15.5 3.73 ;
      RECT  13.01 3.73 15.5 3.735 ;
      RECT  13.005 3.735 15.5 3.74 ;
      RECT  13.0 3.74 15.5 3.745 ;
      RECT  12.995 3.745 15.5 3.75 ;
      RECT  12.99 3.75 15.5 3.755 ;
      RECT  12.985 3.755 15.5 3.76 ;
      RECT  12.98 3.76 15.5 3.765 ;
      RECT  12.975 3.765 15.5 3.77 ;
      RECT  12.97 3.77 15.5 3.775 ;
      RECT  12.965 3.775 15.5 3.78 ;
      RECT  12.96 3.78 15.5 3.785 ;
      RECT  12.955 3.785 15.5 3.79 ;
      RECT  12.95 3.79 15.5 3.795 ;
      RECT  12.945 3.795 15.5 3.8 ;
      RECT  12.94 3.8 15.5 3.805 ;
      RECT  12.935 3.805 15.5 3.81 ;
      RECT  12.93 3.81 15.5 3.815 ;
      RECT  12.925 3.815 15.5 3.82 ;
      RECT  12.92 3.82 15.5 3.825 ;
      RECT  12.915 3.825 15.5 3.83 ;
      RECT  12.91 3.83 15.5 3.835 ;
      RECT  12.905 3.835 15.5 3.84 ;
      RECT  12.9 3.84 15.5 3.845 ;
      RECT  12.895 3.845 15.5 3.85 ;
      RECT  12.89 3.85 15.5 3.855 ;
      RECT  12.885 3.855 15.5 3.86 ;
      RECT  12.88 3.86 15.5 3.865 ;
      RECT  12.875 3.865 15.5 3.87 ;
      RECT  12.87 3.87 15.5 3.875 ;
      RECT  12.865 3.875 15.5 3.88 ;
      RECT  12.86 3.88 15.5 3.885 ;
      RECT  12.855 3.885 15.5 3.89 ;
      RECT  12.85 3.89 15.5 3.895 ;
      RECT  12.845 3.895 15.5 3.9 ;
      RECT  12.84 3.9 15.5 3.905 ;
      RECT  12.835 3.905 15.5 3.91 ;
      RECT  12.83 3.91 15.5 3.915 ;
      RECT  12.825 3.915 13.15 3.92 ;
      RECT  12.82 3.92 13.145 3.925 ;
      RECT  12.815 3.925 13.14 3.93 ;
      RECT  12.81 3.93 13.135 3.935 ;
      RECT  12.805 3.935 13.13 3.94 ;
      RECT  12.8 3.94 13.125 3.945 ;
      RECT  12.795 3.945 13.12 3.95 ;
      RECT  12.79 3.95 13.115 3.955 ;
      RECT  12.785 3.955 13.11 3.96 ;
      RECT  12.78 3.96 13.105 3.965 ;
      RECT  12.775 3.965 13.1 3.97 ;
      RECT  12.77 3.97 13.095 3.975 ;
      RECT  12.765 3.975 13.09 3.98 ;
      RECT  12.76 3.98 13.085 3.985 ;
      RECT  12.755 3.985 13.08 3.99 ;
      RECT  12.75 3.99 13.075 3.995 ;
      RECT  12.745 3.995 13.07 4.0 ;
      RECT  12.74 4.0 13.065 4.005 ;
      RECT  12.735 4.005 13.06 4.01 ;
      RECT  12.73 4.01 13.055 4.015 ;
      RECT  12.725 4.015 13.05 4.02 ;
      RECT  12.72 4.02 13.045 4.025 ;
      RECT  12.715 4.025 13.04 4.03 ;
      RECT  12.71 4.03 13.035 4.035 ;
      RECT  12.705 4.035 13.03 4.04 ;
      RECT  12.7 4.04 13.025 4.045 ;
      RECT  12.695 4.045 13.02 4.05 ;
      RECT  12.69 4.05 13.015 4.055 ;
      RECT  12.685 4.055 13.01 4.06 ;
      RECT  12.68 4.06 13.005 4.065 ;
      RECT  12.675 4.065 13.0 4.07 ;
      RECT  12.67 4.07 12.995 4.075 ;
      RECT  12.665 4.075 12.99 4.08 ;
      RECT  12.66 4.08 12.985 4.085 ;
      RECT  12.655 4.085 12.98 4.09 ;
      RECT  12.65 4.09 12.975 4.095 ;
      RECT  12.645 4.095 12.97 4.1 ;
      RECT  12.64 4.1 12.965 4.105 ;
      RECT  12.635 4.105 12.96 4.11 ;
      RECT  12.63 4.11 12.955 4.115 ;
      RECT  12.625 4.115 12.95 4.12 ;
      RECT  12.62 4.12 12.945 4.125 ;
      RECT  12.615 4.125 12.94 4.13 ;
      RECT  12.61 4.13 12.935 4.135 ;
      RECT  12.605 4.135 12.93 4.14 ;
      RECT  12.6 4.14 12.925 4.145 ;
      RECT  12.595 4.145 12.92 4.15 ;
      RECT  12.59 4.15 12.915 4.155 ;
      RECT  12.585 4.155 12.91 4.16 ;
      RECT  12.58 4.16 12.905 4.165 ;
      RECT  12.575 4.165 12.9 4.17 ;
      RECT  12.57 4.17 12.895 4.175 ;
      RECT  12.565 4.175 12.89 4.18 ;
      RECT  12.56 4.18 12.885 4.185 ;
      RECT  12.555 4.185 12.88 4.19 ;
      RECT  12.55 4.19 12.875 4.195 ;
      RECT  12.545 4.195 12.87 4.2 ;
      RECT  12.54 4.2 12.865 4.205 ;
      RECT  12.535 4.205 12.86 4.21 ;
      RECT  12.53 4.21 12.855 4.215 ;
      RECT  8.75 4.215 12.85 4.22 ;
      RECT  8.75 4.22 12.845 4.225 ;
      RECT  8.75 4.225 12.84 4.23 ;
      RECT  8.75 4.23 12.835 4.235 ;
      RECT  8.75 4.235 12.83 4.24 ;
      RECT  8.75 4.24 12.825 4.245 ;
      RECT  8.75 4.245 12.82 4.25 ;
      RECT  8.75 4.25 12.815 4.255 ;
      RECT  8.75 4.255 12.81 4.26 ;
      RECT  8.75 4.26 12.805 4.265 ;
      RECT  8.75 4.265 12.8 4.27 ;
      RECT  8.75 4.27 12.795 4.275 ;
      RECT  8.75 4.275 12.79 4.28 ;
      RECT  8.75 4.28 12.785 4.285 ;
      RECT  8.75 4.285 12.78 4.29 ;
      RECT  8.75 4.29 12.775 4.295 ;
      RECT  8.75 4.295 12.77 4.3 ;
      RECT  8.75 4.3 12.765 4.305 ;
      RECT  8.75 4.305 12.76 4.31 ;
      RECT  8.75 4.31 12.755 4.315 ;
      RECT  8.75 4.315 12.75 4.32 ;
      RECT  8.75 4.32 12.745 4.325 ;
      RECT  8.75 4.325 12.74 4.33 ;
      RECT  8.75 4.33 12.735 4.335 ;
      RECT  8.75 4.335 12.73 4.34 ;
      RECT  8.75 4.34 12.725 4.345 ;
      RECT  8.75 4.345 12.72 4.35 ;
      RECT  8.75 4.35 12.715 4.355 ;
      RECT  8.75 4.355 12.71 4.36 ;
      RECT  8.75 4.36 12.705 4.365 ;
      RECT  8.75 4.365 12.7 4.37 ;
      RECT  8.75 4.37 12.695 4.375 ;
      RECT  8.75 4.375 12.69 4.38 ;
      RECT  8.75 4.38 12.685 4.385 ;
      RECT  8.75 4.385 12.68 4.39 ;
      RECT  8.75 4.39 12.675 4.395 ;
      RECT  8.75 4.395 12.67 4.4 ;
      RECT  8.75 4.4 12.665 4.405 ;
      RECT  8.75 4.405 12.66 4.41 ;
      RECT  8.75 4.41 12.655 4.415 ;
      RECT  8.75 4.415 12.65 4.42 ;
      RECT  8.75 4.42 12.645 4.425 ;
      RECT  8.75 4.425 12.64 4.43 ;
      RECT  8.75 4.43 12.635 4.435 ;
      RECT  8.75 4.435 12.63 4.44 ;
      RECT  8.75 4.44 12.625 4.445 ;
      RECT  8.75 4.445 8.98 4.48 ;
      RECT  8.44 4.48 8.98 4.71 ;
      RECT  15.745 3.805 18.44 4.035 ;
      RECT  15.745 4.035 15.975 4.16 ;
      RECT  13.525 4.16 15.975 4.39 ;
      RECT  13.525 4.39 13.755 4.48 ;
      RECT  12.92 4.48 13.755 4.71 ;
      RECT  16.205 4.36 16.445 4.365 ;
      RECT  16.205 4.365 17.475 4.595 ;
      RECT  16.205 4.595 16.445 4.62 ;
      RECT  17.245 4.595 17.475 5.0 ;
      RECT  13.985 4.62 16.445 4.85 ;
      RECT  16.205 4.85 16.445 4.855 ;
      RECT  13.985 4.85 14.215 4.98 ;
      RECT  12.205 4.87 12.435 4.98 ;
      RECT  12.205 4.98 14.215 5.21 ;
      RECT  17.19 5.0 17.53 5.23 ;
      RECT  4.365 4.215 7.24 4.445 ;
      RECT  4.365 4.445 4.595 4.525 ;
      RECT  3.19 4.525 4.595 4.755 ;
      RECT  9.21 4.675 10.755 4.905 ;
      RECT  9.21 4.905 9.44 5.0 ;
      RECT  10.525 4.905 10.755 5.0 ;
      RECT  8.23 5.0 9.44 5.23 ;
      RECT  10.525 5.0 11.93 5.23 ;
      LAYER METAL2 ;
      RECT  8.77 2.66 10.83 2.94 ;
      RECT  7.115 3.22 9.635 3.5 ;
      LAYER VIA12 ;
      RECT  8.83 2.67 9.09 2.93 ;
      RECT  10.51 2.67 10.77 2.93 ;
      RECT  7.175 3.23 7.435 3.49 ;
      RECT  9.23 3.23 9.49 3.49 ;
  END
END MDN_FSDNRB_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNRB_1
#      Description : D-Flip Flop w/scan, neg-edge triggered, lo-async-clear
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNRB_1
  CLASS CORE ;
  FOREIGN MDN_FSDNRB_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.405 2.1 10.195 2.38 ;
      RECT  9.405 2.38 9.635 2.69 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  20.3 1.565 21.395 1.795 ;
      RECT  21.165 1.795 21.395 3.245 ;
      RECT  20.34 3.245 21.395 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  21.725 1.565 22.22 1.795 ;
      RECT  21.725 1.795 21.955 3.245 ;
      RECT  21.725 3.245 22.22 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END QN
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  16.125 4.635 17.475 4.865 ;
      RECT  16.125 4.865 16.355 4.925 ;
      RECT  17.245 4.865 17.475 5.0 ;
      RECT  13.325 4.925 16.355 5.0 ;
      RECT  9.505 4.41 12.94 4.64 ;
      RECT  9.505 4.64 9.735 5.0 ;
      RECT  12.71 4.64 12.94 5.0 ;
      RECT  3.75 5.0 9.735 5.23 ;
      RECT  12.71 5.0 16.355 5.155 ;
      RECT  17.245 5.0 18.65 5.23 ;
      RECT  18.34 4.365 18.62 5.0 ;
      RECT  12.71 5.155 13.555 5.23 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.63 5.095 16.97 5.46 ;
      RECT  16.24 5.46 17.36 5.74 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.73 ;
      RECT  18.365 -0.14 19.04 0.14 ;
      RECT  18.365 0.14 18.595 1.005 ;
      RECT  18.1 1.005 18.595 1.235 ;
      RECT  16.24 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.6 ;
      RECT  9.965 -0.14 12.995 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  12.765 0.14 12.995 1.005 ;
      RECT  12.765 1.005 13.26 1.235 ;
      RECT  6.045 -0.14 6.72 0.14 ;
      RECT  6.045 0.14 6.275 0.89 ;
      RECT  6.045 0.89 6.54 1.12 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 10.81 0.445 ;
      RECT  10.47 0.445 12.435 0.675 ;
      RECT  12.205 0.675 12.435 1.525 ;
      RECT  12.205 1.525 14.115 1.655 ;
      RECT  12.205 1.655 14.89 1.755 ;
      RECT  13.885 1.755 14.89 1.885 ;
      RECT  14.66 1.885 14.89 2.335 ;
      RECT  14.66 2.335 15.29 2.565 ;
      RECT  21.67 0.37 22.01 0.6 ;
      RECT  21.67 0.6 21.9 1.005 ;
      RECT  18.925 0.37 20.835 0.6 ;
      RECT  20.605 0.6 20.835 1.005 ;
      RECT  18.925 0.6 19.155 1.565 ;
      RECT  20.605 1.005 21.9 1.235 ;
      RECT  14.385 1.005 15.795 1.235 ;
      RECT  15.565 1.235 15.795 1.29 ;
      RECT  15.565 1.29 17.05 1.52 ;
      RECT  16.82 1.52 17.05 1.565 ;
      RECT  16.82 1.565 19.155 1.795 ;
      RECT  16.82 1.795 17.05 3.715 ;
      RECT  14.39 3.715 17.05 3.945 ;
      RECT  3.19 0.445 4.595 0.675 ;
      RECT  4.365 0.675 4.595 1.005 ;
      RECT  4.365 1.005 5.0 1.235 ;
      RECT  13.675 0.445 16.355 0.675 ;
      RECT  16.125 0.675 16.355 0.83 ;
      RECT  13.675 0.675 13.905 1.29 ;
      RECT  16.125 0.83 17.74 1.06 ;
      RECT  17.4 1.06 17.74 1.12 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  8.44 1.005 11.72 1.235 ;
      RECT  19.485 1.005 19.98 1.235 ;
      RECT  19.485 1.235 19.715 2.125 ;
      RECT  17.28 2.125 20.835 2.355 ;
      RECT  17.28 2.355 17.51 2.685 ;
      RECT  20.605 2.355 20.835 2.69 ;
      RECT  18.365 2.355 18.595 3.245 ;
      RECT  19.485 2.355 19.715 3.245 ;
      RECT  18.1 3.245 18.595 3.475 ;
      RECT  19.485 3.245 19.98 3.475 ;
      RECT  6.045 1.47 7.24 1.565 ;
      RECT  3.96 1.565 7.24 1.7 ;
      RECT  3.96 1.7 6.275 1.795 ;
      RECT  1.72 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 3.245 ;
      RECT  1.72 3.245 6.275 3.475 ;
      RECT  6.045 2.35 6.275 3.245 ;
      RECT  8.845 1.565 9.48 1.795 ;
      RECT  8.845 1.795 9.075 2.335 ;
      RECT  8.23 2.335 9.075 2.565 ;
      RECT  8.845 2.565 9.075 3.03 ;
      RECT  8.845 3.03 10.755 3.26 ;
      RECT  10.525 2.35 10.755 3.03 ;
      RECT  10.68 1.565 11.315 1.795 ;
      RECT  11.085 1.795 11.315 1.985 ;
      RECT  11.085 1.985 13.555 2.215 ;
      RECT  13.325 2.215 13.555 2.335 ;
      RECT  11.085 2.215 11.315 3.49 ;
      RECT  13.325 2.335 14.17 2.565 ;
      RECT  7.165 2.39 7.395 2.795 ;
      RECT  7.165 2.795 8.515 3.025 ;
      RECT  8.285 3.025 8.515 3.49 ;
      RECT  8.285 3.49 11.315 3.72 ;
      RECT  7.725 1.695 7.955 1.93 ;
      RECT  6.605 1.93 7.955 2.16 ;
      RECT  6.605 2.16 6.835 3.22 ;
      RECT  6.605 3.22 6.985 3.255 ;
      RECT  6.605 3.255 8.01 3.485 ;
      RECT  6.605 3.485 6.985 3.5 ;
      RECT  15.16 1.75 16.59 1.98 ;
      RECT  16.36 1.98 16.59 3.255 ;
      RECT  13.62 3.255 16.59 3.485 ;
      RECT  13.62 3.485 13.85 3.805 ;
      RECT  11.815 2.445 12.435 2.675 ;
      RECT  12.205 2.675 12.435 3.805 ;
      RECT  12.205 3.805 13.85 4.035 ;
      RECT  15.9 2.39 16.13 2.795 ;
      RECT  13.03 2.795 16.13 3.025 ;
      RECT  13.03 3.025 13.26 3.22 ;
      RECT  12.665 3.22 13.26 3.5 ;
      RECT  5.42 3.805 7.955 4.025 ;
      RECT  5.42 4.025 8.78 4.035 ;
      RECT  7.725 4.035 8.78 4.255 ;
      RECT  2.41 3.805 5.0 4.035 ;
      RECT  9.035 3.95 11.72 4.18 ;
      RECT  9.035 4.18 9.265 4.485 ;
      RECT  6.955 4.31 7.185 4.485 ;
      RECT  6.955 4.485 9.265 4.715 ;
      RECT  15.16 4.175 17.74 4.405 ;
      RECT  0.14 4.365 6.54 4.595 ;
      RECT  1.51 5.0 2.97 5.23 ;
      LAYER METAL2 ;
      RECT  6.605 3.22 13.045 3.5 ;
      LAYER VIA12 ;
      RECT  6.665 3.23 6.925 3.49 ;
      RECT  12.725 3.23 12.985 3.49 ;
  END
END MDN_FSDNRB_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNRB_2
#      Description : D-Flip Flop w/scan, neg-edge triggered, lo-async-clear
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNRB_2
  CLASS CORE ;
  FOREIGN MDN_FSDNRB_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 24.64 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.405 2.1 10.195 2.38 ;
      RECT  9.405 2.38 9.635 2.69 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  20.34 1.565 22.22 1.795 ;
      RECT  21.165 1.795 21.395 3.245 ;
      RECT  20.34 3.245 22.22 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  22.58 1.565 24.46 1.795 ;
      RECT  23.405 1.795 23.635 3.245 ;
      RECT  22.58 3.245 24.46 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END QN
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  16.125 4.67 17.475 4.9 ;
      RECT  16.125 4.9 16.355 4.925 ;
      RECT  17.245 4.9 17.475 5.0 ;
      RECT  13.325 4.925 16.355 5.0 ;
      RECT  9.505 4.515 12.92 4.745 ;
      RECT  9.505 4.745 9.735 4.925 ;
      RECT  12.69 4.745 12.92 5.0 ;
      RECT  4.365 4.925 9.735 5.0 ;
      RECT  3.75 5.0 9.735 5.155 ;
      RECT  12.69 5.0 16.355 5.155 ;
      RECT  17.245 5.0 18.65 5.23 ;
      RECT  18.34 4.365 18.62 5.0 ;
      RECT  3.75 5.155 4.595 5.23 ;
      RECT  12.69 5.155 13.555 5.23 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 2.94 2.355 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.81 5.74 ;
      RECT  21.165 4.87 21.395 5.46 ;
      RECT  21.165 5.46 21.84 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.63 5.135 16.97 5.46 ;
      RECT  16.24 5.46 17.36 5.74 ;
      RECT  9.965 4.975 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.975 12.435 5.46 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 24.64 5.74 ;
      LAYER VIA12 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  24.23 5.47 24.49 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 -0.14 24.81 0.14 ;
      RECT  23.405 0.14 23.635 0.73 ;
      RECT  21.165 -0.14 21.84 0.14 ;
      RECT  21.165 0.14 21.395 0.73 ;
      RECT  18.365 -0.14 19.04 0.14 ;
      RECT  18.365 0.14 18.595 1.005 ;
      RECT  18.1 1.005 18.595 1.235 ;
      RECT  16.24 -0.14 17.36 0.14 ;
      RECT  16.63 0.14 16.97 0.465 ;
      RECT  9.965 -0.14 12.995 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  12.765 0.14 12.995 1.005 ;
      RECT  12.765 1.005 13.26 1.235 ;
      RECT  6.045 -0.14 6.72 0.14 ;
      RECT  6.045 0.14 6.275 0.89 ;
      RECT  6.045 0.89 6.54 1.12 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 24.64 0.14 ;
      LAYER VIA12 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 12.435 0.6 ;
      RECT  12.205 0.6 12.435 1.525 ;
      RECT  12.205 1.525 14.13 1.635 ;
      RECT  12.205 1.635 14.675 1.755 ;
      RECT  13.9 1.755 14.675 1.865 ;
      RECT  14.445 1.865 14.675 2.335 ;
      RECT  14.445 2.335 15.29 2.565 ;
      RECT  23.91 0.37 24.25 0.6 ;
      RECT  23.91 0.6 24.14 1.005 ;
      RECT  22.79 0.37 23.13 0.6 ;
      RECT  22.79 0.6 23.02 1.005 ;
      RECT  19.43 0.37 19.77 0.6 ;
      RECT  19.43 0.6 19.66 1.005 ;
      RECT  18.925 1.005 24.14 1.235 ;
      RECT  18.925 1.235 19.155 1.565 ;
      RECT  14.39 1.155 17.05 1.385 ;
      RECT  16.82 1.385 17.05 1.565 ;
      RECT  16.82 1.565 19.155 1.795 ;
      RECT  16.82 1.795 17.05 3.715 ;
      RECT  14.39 3.715 17.05 3.945 ;
      RECT  13.675 0.695 17.685 0.925 ;
      RECT  13.675 0.925 13.905 1.29 ;
      RECT  17.455 0.925 17.685 1.29 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.19 1.005 5.0 1.235 ;
      RECT  8.44 1.005 11.72 1.235 ;
      RECT  6.045 1.465 7.24 1.565 ;
      RECT  3.96 1.565 7.24 1.695 ;
      RECT  3.96 1.695 6.275 1.795 ;
      RECT  1.72 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 3.245 ;
      RECT  1.72 3.245 6.275 3.475 ;
      RECT  6.045 2.35 6.275 3.245 ;
      RECT  8.845 1.565 9.48 1.795 ;
      RECT  8.845 1.795 9.075 2.335 ;
      RECT  8.23 2.335 9.075 2.565 ;
      RECT  8.845 2.565 9.075 3.03 ;
      RECT  8.845 3.03 10.755 3.26 ;
      RECT  10.525 2.35 10.755 3.03 ;
      RECT  10.68 1.565 11.315 1.795 ;
      RECT  11.085 1.795 11.315 1.985 ;
      RECT  11.085 1.985 13.65 2.215 ;
      RECT  13.42 2.215 13.65 2.335 ;
      RECT  11.085 2.215 11.315 3.545 ;
      RECT  13.42 2.335 14.17 2.565 ;
      RECT  7.165 2.39 7.395 2.795 ;
      RECT  7.165 2.795 8.515 3.025 ;
      RECT  8.285 3.025 8.515 3.545 ;
      RECT  8.285 3.545 11.315 3.775 ;
      RECT  19.485 1.565 19.98 1.795 ;
      RECT  19.485 1.795 19.715 2.125 ;
      RECT  17.28 2.125 20.835 2.355 ;
      RECT  17.28 2.355 17.51 2.69 ;
      RECT  20.605 2.355 20.835 2.69 ;
      RECT  18.365 2.355 18.595 3.245 ;
      RECT  19.485 2.355 19.715 3.245 ;
      RECT  18.1 3.245 18.595 3.475 ;
      RECT  19.485 3.245 19.98 3.475 ;
      RECT  15.16 1.615 16.59 1.845 ;
      RECT  16.36 1.845 16.59 3.255 ;
      RECT  13.62 3.255 16.59 3.485 ;
      RECT  13.62 3.485 13.85 3.805 ;
      RECT  11.59 2.445 12.435 2.675 ;
      RECT  12.205 2.675 12.435 3.805 ;
      RECT  12.205 3.805 13.85 4.035 ;
      RECT  7.725 1.695 7.955 1.93 ;
      RECT  6.605 1.93 7.955 2.16 ;
      RECT  6.605 2.16 6.835 3.22 ;
      RECT  6.605 3.22 6.985 3.255 ;
      RECT  6.605 3.255 8.01 3.485 ;
      RECT  6.605 3.485 6.985 3.5 ;
      RECT  15.9 2.35 16.13 2.795 ;
      RECT  13.03 2.795 16.13 3.025 ;
      RECT  13.03 3.025 13.26 3.22 ;
      RECT  12.69 3.22 13.26 3.5 ;
      RECT  5.43 3.805 7.395 4.005 ;
      RECT  5.43 4.005 8.78 4.035 ;
      RECT  7.165 4.035 8.78 4.235 ;
      RECT  2.42 3.805 5.0 4.035 ;
      RECT  9.035 4.045 11.72 4.275 ;
      RECT  9.035 4.275 9.265 4.465 ;
      RECT  6.9 4.465 9.265 4.695 ;
      RECT  15.16 4.175 17.74 4.405 ;
      RECT  0.18 4.365 6.54 4.595 ;
      RECT  20.66 4.365 21.9 4.595 ;
      RECT  20.66 4.595 20.89 5.0 ;
      RECT  21.67 4.595 21.9 5.0 ;
      RECT  20.55 5.0 20.89 5.23 ;
      RECT  21.67 5.0 22.01 5.23 ;
      LAYER METAL2 ;
      RECT  6.605 3.22 13.07 3.5 ;
      LAYER VIA12 ;
      RECT  6.665 3.23 6.925 3.49 ;
      RECT  12.75 3.23 13.01 3.49 ;
  END
END MDN_FSDNRB_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNRBQ_F_1
#      Description : D-Flip Flop w/scan, neg-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNRBQ_F_1
  CLASS CORE ;
  FOREIGN MDN_FSDNRBQ_F_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  21.725 1.565 22.22 1.795 ;
      RECT  21.725 1.795 21.955 3.245 ;
      RECT  21.725 3.245 22.22 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 2.445 13.05 2.675 ;
      RECT  12.205 2.675 12.435 3.245 ;
      RECT  10.525 3.245 12.435 3.475 ;
      RECT  10.525 3.475 10.755 3.49 ;
      RECT  12.205 3.475 12.435 3.98 ;
      RECT  8.26 2.125 8.54 3.49 ;
      RECT  8.26 3.49 10.755 3.72 ;
      RECT  12.205 3.98 15.595 4.21 ;
      RECT  15.365 4.21 15.595 4.54 ;
      RECT  15.365 4.54 19.64 4.77 ;
      RECT  19.41 4.77 19.64 5.0 ;
      RECT  19.41 5.0 19.77 5.23 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.87 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 5.08 19.155 5.46 ;
      RECT  18.925 5.46 20.16 5.74 ;
      RECT  12.205 4.93 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 4.93 14.675 5.46 ;
      RECT  7.725 4.93 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.19 5.135 3.53 5.46 ;
      RECT  2.8 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  19.6 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  20.045 0.14 20.275 1.005 ;
      RECT  19.64 1.005 20.275 1.235 ;
      RECT  12.765 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.765 0.14 12.995 1.005 ;
      RECT  12.765 1.005 13.26 1.235 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.6 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  20.31 -0.13 20.57 0.13 ;
      RECT  20.87 -0.13 21.13 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.5 0.37 1.85 0.6 ;
      RECT  1.5 0.6 1.73 1.005 ;
      RECT  0.18 1.005 1.73 1.235 ;
      RECT  2.63 0.37 7.45 0.6 ;
      RECT  9.35 0.37 10.195 0.6 ;
      RECT  9.965 0.6 10.195 0.98 ;
      RECT  9.89 0.98 10.27 1.26 ;
      RECT  11.59 0.37 12.435 0.6 ;
      RECT  12.205 0.6 12.435 1.525 ;
      RECT  12.205 1.525 14.675 1.755 ;
      RECT  14.445 1.755 14.675 2.405 ;
      RECT  14.445 2.405 15.29 2.635 ;
      RECT  14.445 2.635 14.675 3.52 ;
      RECT  13.62 3.52 14.675 3.75 ;
      RECT  16.685 0.37 17.53 0.6 ;
      RECT  16.685 0.6 16.915 1.005 ;
      RECT  13.81 0.98 14.19 1.005 ;
      RECT  13.81 1.005 16.915 1.235 ;
      RECT  13.81 1.235 14.19 1.26 ;
      RECT  18.31 0.37 19.155 0.6 ;
      RECT  18.925 0.6 19.155 1.565 ;
      RECT  18.925 1.565 20.68 1.795 ;
      RECT  18.925 1.795 19.155 3.16 ;
      RECT  18.925 3.16 20.68 3.39 ;
      RECT  2.61 0.98 2.99 1.005 ;
      RECT  1.96 1.005 2.99 1.235 ;
      RECT  2.61 1.235 2.99 1.26 ;
      RECT  1.96 1.235 2.19 1.565 ;
      RECT  1.565 1.565 2.19 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 2.06 4.035 ;
      RECT  4.925 0.83 9.425 1.005 ;
      RECT  3.245 1.005 9.425 1.06 ;
      RECT  3.245 1.06 5.155 1.235 ;
      RECT  9.195 1.06 9.425 1.29 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  2.42 1.565 3.475 1.795 ;
      RECT  10.68 1.005 11.72 1.235 ;
      RECT  17.4 1.005 18.44 1.235 ;
      RECT  6.31 1.29 8.515 1.52 ;
      RECT  6.31 1.52 6.54 1.565 ;
      RECT  8.285 1.52 8.515 1.565 ;
      RECT  3.96 1.565 6.54 1.795 ;
      RECT  8.285 1.565 8.78 1.795 ;
      RECT  15.16 1.565 16.2 1.795 ;
      RECT  15.565 1.795 15.795 2.685 ;
      RECT  15.565 2.685 17.475 2.915 ;
      RECT  17.245 2.915 17.475 3.115 ;
      RECT  15.565 2.915 15.795 3.245 ;
      RECT  17.245 3.115 17.74 3.345 ;
      RECT  15.16 3.245 15.795 3.475 ;
      RECT  6.9 1.75 7.395 1.98 ;
      RECT  7.165 1.98 7.395 2.42 ;
      RECT  5.99 2.42 7.395 2.65 ;
      RECT  7.165 2.65 7.395 3.245 ;
      RECT  6.9 3.245 7.395 3.475 ;
      RECT  9.965 1.51 10.195 1.985 ;
      RECT  9.965 1.985 14.115 2.215 ;
      RECT  9.965 2.215 10.195 3.03 ;
      RECT  13.885 2.215 14.115 3.06 ;
      RECT  9.91 3.03 10.25 3.26 ;
      RECT  12.92 3.06 14.115 3.29 ;
      RECT  16.685 1.51 16.915 2.125 ;
      RECT  16.685 2.125 18.595 2.355 ;
      RECT  18.365 2.355 18.595 3.62 ;
      RECT  16.63 3.62 20.78 3.85 ;
      RECT  20.55 3.85 20.78 4.365 ;
      RECT  20.55 4.365 21.9 4.595 ;
      RECT  20.55 4.595 20.78 5.0 ;
      RECT  21.67 4.595 21.9 5.0 ;
      RECT  20.55 5.0 20.89 5.23 ;
      RECT  21.67 5.0 22.01 5.23 ;
      RECT  5.43 3.805 7.965 3.95 ;
      RECT  5.43 3.95 11.02 4.035 ;
      RECT  7.705 4.035 11.02 4.18 ;
      RECT  2.42 3.755 5.0 3.985 ;
      RECT  2.42 3.985 2.76 4.035 ;
      RECT  11.285 3.805 11.72 4.035 ;
      RECT  11.285 4.035 11.515 4.41 ;
      RECT  9.14 4.41 11.515 4.64 ;
      RECT  15.86 4.08 19.98 4.31 ;
      RECT  3.96 4.215 4.595 4.365 ;
      RECT  3.96 4.365 6.54 4.445 ;
      RECT  4.365 4.445 6.54 4.595 ;
      RECT  11.745 4.44 15.135 4.67 ;
      RECT  11.745 4.67 11.975 5.0 ;
      RECT  14.905 4.67 15.135 5.0 ;
      RECT  7.16 4.47 8.77 4.7 ;
      RECT  7.16 4.7 7.39 4.925 ;
      RECT  8.54 4.7 8.77 5.0 ;
      RECT  0.18 4.365 3.475 4.595 ;
      RECT  3.245 4.595 3.475 4.675 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  3.245 4.675 4.035 4.905 ;
      RECT  3.805 4.905 4.035 4.925 ;
      RECT  3.805 4.925 7.39 5.155 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  8.54 5.0 11.975 5.23 ;
      RECT  14.905 5.0 16.41 5.23 ;
      LAYER METAL2 ;
      RECT  2.61 0.98 14.19 1.26 ;
      LAYER VIA12 ;
      RECT  2.67 0.99 2.93 1.25 ;
      RECT  9.95 0.99 10.21 1.25 ;
      RECT  13.87 0.99 14.13 1.25 ;
  END
END MDN_FSDNRBQ_F_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNRBQ_F_2
#      Description : D-Flip Flop w/scan, neg-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNRBQ_F_2
  CLASS CORE ;
  FOREIGN MDN_FSDNRBQ_F_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 24.64 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  21.88 1.565 22.92 1.795 ;
      RECT  22.285 1.795 22.515 3.245 ;
      RECT  21.88 3.245 22.92 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 2.445 13.05 2.675 ;
      RECT  12.205 2.675 12.435 3.245 ;
      RECT  10.525 3.245 12.435 3.475 ;
      RECT  10.525 3.475 10.755 3.49 ;
      RECT  12.205 3.475 12.435 4.06 ;
      RECT  8.26 2.125 8.54 3.49 ;
      RECT  8.26 3.49 10.755 3.72 ;
      RECT  12.205 4.06 12.995 4.165 ;
      RECT  12.205 4.165 15.65 4.29 ;
      RECT  12.765 4.29 15.65 4.395 ;
      RECT  15.42 4.395 15.65 4.54 ;
      RECT  15.42 4.54 19.64 4.77 ;
      RECT  19.41 4.77 19.64 5.0 ;
      RECT  19.41 5.0 19.77 5.23 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.81 5.74 ;
      RECT  21.165 4.87 21.395 5.46 ;
      RECT  21.165 5.46 22.4 5.74 ;
      RECT  18.925 5.0 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  12.15 5.135 12.49 5.46 ;
      RECT  11.76 5.46 15.12 5.74 ;
      RECT  14.39 5.135 14.73 5.46 ;
      RECT  7.725 4.93 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.19 5.135 3.53 5.46 ;
      RECT  2.8 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 24.64 5.74 ;
      LAYER VIA12 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  24.23 5.47 24.49 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 -0.14 24.81 0.14 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  19.6 -0.14 21.395 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  20.045 0.14 20.275 1.005 ;
      RECT  19.64 1.005 20.275 1.235 ;
      RECT  12.32 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.765 0.14 12.995 1.005 ;
      RECT  12.765 1.005 13.26 1.235 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.6 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 24.64 0.14 ;
      LAYER VIA12 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  20.31 -0.13 20.57 0.13 ;
      RECT  20.87 -0.13 21.13 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  17.19 0.37 17.53 0.44 ;
      RECT  15.005 0.44 17.53 0.67 ;
      RECT  15.005 0.67 15.235 1.005 ;
      RECT  13.81 0.98 14.19 1.005 ;
      RECT  13.81 1.005 15.235 1.235 ;
      RECT  13.81 1.235 14.19 1.26 ;
      RECT  1.465 0.37 1.85 0.6 ;
      RECT  1.465 0.6 1.695 1.005 ;
      RECT  0.18 1.005 1.695 1.235 ;
      RECT  2.63 0.37 7.45 0.6 ;
      RECT  9.35 0.37 10.195 0.6 ;
      RECT  9.965 0.6 10.195 0.98 ;
      RECT  9.89 0.98 10.27 1.26 ;
      RECT  11.59 0.37 12.435 0.6 ;
      RECT  12.205 0.6 12.435 1.525 ;
      RECT  12.205 1.525 14.675 1.755 ;
      RECT  14.445 1.755 14.675 2.41 ;
      RECT  14.445 2.41 15.29 2.64 ;
      RECT  14.445 2.64 14.675 3.705 ;
      RECT  13.62 3.705 14.675 3.935 ;
      RECT  18.31 0.37 19.155 0.6 ;
      RECT  18.925 0.6 19.155 1.565 ;
      RECT  18.925 1.565 20.68 1.795 ;
      RECT  18.925 1.795 19.155 3.16 ;
      RECT  18.925 3.16 20.68 3.39 ;
      RECT  2.61 0.98 2.99 1.005 ;
      RECT  1.94 1.005 2.99 1.235 ;
      RECT  2.61 1.235 2.99 1.26 ;
      RECT  1.94 1.235 2.17 1.565 ;
      RECT  1.565 1.565 2.17 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 2.06 4.035 ;
      RECT  4.92 0.83 9.425 1.005 ;
      RECT  3.24 1.005 9.425 1.06 ;
      RECT  3.24 1.06 5.155 1.235 ;
      RECT  9.195 1.06 9.425 1.29 ;
      RECT  3.24 1.235 3.47 1.565 ;
      RECT  2.42 1.565 3.47 1.795 ;
      RECT  10.68 1.005 11.72 1.235 ;
      RECT  17.4 1.005 18.44 1.235 ;
      RECT  6.31 1.29 8.515 1.52 ;
      RECT  6.31 1.52 6.54 1.565 ;
      RECT  8.285 1.52 8.515 1.565 ;
      RECT  3.96 1.565 6.54 1.795 ;
      RECT  8.285 1.565 8.78 1.795 ;
      RECT  15.16 1.565 16.355 1.795 ;
      RECT  16.125 1.795 16.355 3.03 ;
      RECT  16.125 3.03 17.74 3.245 ;
      RECT  15.16 3.245 17.74 3.26 ;
      RECT  15.16 3.26 16.355 3.475 ;
      RECT  6.9 1.75 7.24 1.98 ;
      RECT  6.9 1.98 7.13 2.405 ;
      RECT  5.99 2.405 7.13 2.635 ;
      RECT  6.9 2.635 7.13 3.245 ;
      RECT  6.9 3.245 7.24 3.475 ;
      RECT  9.965 1.51 10.195 1.985 ;
      RECT  9.965 1.985 14.115 2.215 ;
      RECT  9.965 2.215 10.195 3.03 ;
      RECT  13.885 2.215 14.115 3.245 ;
      RECT  9.91 3.03 10.25 3.26 ;
      RECT  12.92 3.245 14.115 3.475 ;
      RECT  16.685 1.51 16.915 2.125 ;
      RECT  16.685 2.125 18.595 2.355 ;
      RECT  18.365 2.355 18.595 3.62 ;
      RECT  16.63 3.62 20.89 3.85 ;
      RECT  20.66 3.85 20.89 4.37 ;
      RECT  20.66 4.37 21.9 4.6 ;
      RECT  20.66 4.6 20.89 5.0 ;
      RECT  21.67 4.6 21.9 5.0 ;
      RECT  20.55 5.0 20.89 5.23 ;
      RECT  21.67 5.0 23.13 5.23 ;
      RECT  3.5 3.75 4.945 3.805 ;
      RECT  2.42 3.805 4.945 3.98 ;
      RECT  2.42 3.98 3.73 4.035 ;
      RECT  4.715 3.98 4.945 4.09 ;
      RECT  5.43 3.805 7.925 3.95 ;
      RECT  5.43 3.95 11.02 4.035 ;
      RECT  7.705 4.035 11.02 4.18 ;
      RECT  11.25 3.805 11.72 4.035 ;
      RECT  11.25 4.035 11.48 4.33 ;
      RECT  11.245 4.33 11.48 4.335 ;
      RECT  11.24 4.335 11.48 4.34 ;
      RECT  11.235 4.34 11.48 4.345 ;
      RECT  11.23 4.345 11.48 4.35 ;
      RECT  11.225 4.35 11.48 4.355 ;
      RECT  11.22 4.355 11.48 4.36 ;
      RECT  11.215 4.36 11.48 4.365 ;
      RECT  11.21 4.365 11.48 4.37 ;
      RECT  11.205 4.37 11.48 4.375 ;
      RECT  11.2 4.375 11.48 4.38 ;
      RECT  11.195 4.38 11.48 4.385 ;
      RECT  11.19 4.385 11.48 4.39 ;
      RECT  11.185 4.39 11.48 4.395 ;
      RECT  11.18 4.395 11.48 4.4 ;
      RECT  11.175 4.4 11.48 4.405 ;
      RECT  11.17 4.405 11.48 4.41 ;
      RECT  9.14 4.41 11.48 4.425 ;
      RECT  9.14 4.425 11.475 4.43 ;
      RECT  9.14 4.43 11.47 4.435 ;
      RECT  9.14 4.435 11.465 4.44 ;
      RECT  9.14 4.44 11.46 4.445 ;
      RECT  9.14 4.445 11.455 4.45 ;
      RECT  9.14 4.45 11.45 4.455 ;
      RECT  9.14 4.455 11.445 4.46 ;
      RECT  9.14 4.46 11.44 4.465 ;
      RECT  9.14 4.465 11.435 4.47 ;
      RECT  9.14 4.47 11.43 4.475 ;
      RECT  9.14 4.475 11.425 4.48 ;
      RECT  9.14 4.48 11.42 4.485 ;
      RECT  9.14 4.485 11.415 4.49 ;
      RECT  9.14 4.49 11.41 4.495 ;
      RECT  9.14 4.495 11.405 4.5 ;
      RECT  9.14 4.5 11.4 4.505 ;
      RECT  9.14 4.505 11.395 4.51 ;
      RECT  9.14 4.51 11.39 4.515 ;
      RECT  9.14 4.515 11.385 4.52 ;
      RECT  9.14 4.52 11.38 4.525 ;
      RECT  9.14 4.525 11.375 4.53 ;
      RECT  9.14 4.53 11.37 4.535 ;
      RECT  9.14 4.535 11.365 4.54 ;
      RECT  9.14 4.54 11.36 4.545 ;
      RECT  9.14 4.545 11.355 4.55 ;
      RECT  9.14 4.55 11.35 4.555 ;
      RECT  9.14 4.555 11.345 4.56 ;
      RECT  9.14 4.56 11.34 4.565 ;
      RECT  9.14 4.565 11.335 4.57 ;
      RECT  9.14 4.57 11.33 4.575 ;
      RECT  9.14 4.575 11.325 4.58 ;
      RECT  9.14 4.58 11.32 4.585 ;
      RECT  9.14 4.585 11.315 4.59 ;
      RECT  9.14 4.59 11.31 4.595 ;
      RECT  9.14 4.595 11.305 4.6 ;
      RECT  9.14 4.6 11.3 4.605 ;
      RECT  9.14 4.605 11.295 4.61 ;
      RECT  9.14 4.61 11.29 4.615 ;
      RECT  9.14 4.615 11.285 4.62 ;
      RECT  9.14 4.62 11.28 4.625 ;
      RECT  9.14 4.625 11.275 4.63 ;
      RECT  9.14 4.63 11.27 4.635 ;
      RECT  9.14 4.635 11.265 4.64 ;
      RECT  15.86 3.805 16.355 4.035 ;
      RECT  16.125 4.035 16.355 4.08 ;
      RECT  16.125 4.08 19.98 4.31 ;
      RECT  3.96 4.215 4.49 4.365 ;
      RECT  3.96 4.365 6.54 4.445 ;
      RECT  4.26 4.445 6.54 4.595 ;
      RECT  11.69 4.675 15.19 4.905 ;
      RECT  11.69 4.905 11.92 5.0 ;
      RECT  14.96 4.905 15.19 5.0 ;
      RECT  7.165 4.47 8.515 4.7 ;
      RECT  7.165 4.7 7.395 4.925 ;
      RECT  8.285 4.7 8.515 5.0 ;
      RECT  0.18 4.365 2.915 4.595 ;
      RECT  2.685 4.595 2.915 4.675 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  2.685 4.675 4.035 4.905 ;
      RECT  3.805 4.905 4.035 4.925 ;
      RECT  3.805 4.925 7.395 5.155 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  8.285 5.0 11.92 5.23 ;
      RECT  14.96 5.0 16.42 5.23 ;
      LAYER METAL2 ;
      RECT  2.61 0.98 14.19 1.26 ;
      LAYER VIA12 ;
      RECT  2.67 0.99 2.93 1.25 ;
      RECT  9.95 0.99 10.21 1.25 ;
      RECT  13.87 0.99 14.13 1.25 ;
  END
END MDN_FSDNRBQ_F_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNRBQ_F_4
#      Description : D-Flip Flop w/scan, neg-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNRBQ_F_4
  CLASS CORE ;
  FOREIGN MDN_FSDNRBQ_F_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 26.88 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  21.88 1.565 25.16 1.795 ;
      RECT  23.405 1.795 23.635 3.245 ;
      RECT  21.88 3.245 25.16 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 2.445 13.05 2.675 ;
      RECT  12.205 2.675 12.435 3.245 ;
      RECT  11.085 3.245 12.435 3.475 ;
      RECT  11.085 3.475 11.315 3.49 ;
      RECT  12.205 3.475 12.435 3.95 ;
      RECT  8.26 2.125 8.54 2.915 ;
      RECT  8.285 2.915 8.515 3.49 ;
      RECT  8.285 3.49 11.315 3.72 ;
      RECT  12.205 3.95 15.595 4.18 ;
      RECT  15.365 4.18 15.595 4.54 ;
      RECT  15.365 4.54 19.64 4.77 ;
      RECT  19.41 4.77 19.64 5.0 ;
      RECT  19.41 5.0 19.77 5.23 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.645 5.46 27.05 5.74 ;
      RECT  23.405 4.87 23.635 5.46 ;
      RECT  22.96 5.46 23.635 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  20.72 5.46 21.395 5.74 ;
      RECT  18.925 5.0 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  12.205 5.08 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 5.08 14.675 5.46 ;
      RECT  7.725 4.93 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.19 5.135 3.53 5.46 ;
      RECT  2.8 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 26.88 5.74 ;
      LAYER VIA12 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 -0.14 27.05 0.14 ;
      RECT  25.645 0.14 25.875 0.7 ;
      RECT  22.96 -0.14 23.635 0.14 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  21.165 -0.14 21.84 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  19.04 -0.14 19.715 0.14 ;
      RECT  19.485 0.14 19.715 1.005 ;
      RECT  19.485 1.005 19.98 1.235 ;
      RECT  12.765 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.765 0.14 12.995 1.005 ;
      RECT  12.765 1.005 13.26 1.235 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.6 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 26.88 0.14 ;
      LAYER VIA12 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  23.11 -0.13 23.37 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  2.63 0.37 2.97 0.445 ;
      RECT  2.63 0.445 7.45 0.6 ;
      RECT  5.49 0.37 7.45 0.445 ;
      RECT  2.63 0.6 5.715 0.675 ;
      RECT  1.5 0.37 1.85 0.6 ;
      RECT  1.5 0.6 1.73 1.005 ;
      RECT  0.18 1.005 1.73 1.235 ;
      RECT  9.35 0.37 10.19 0.6 ;
      RECT  9.96 0.6 10.19 0.98 ;
      RECT  9.89 0.98 10.27 1.26 ;
      RECT  11.59 0.37 12.435 0.6 ;
      RECT  12.205 0.6 12.435 1.525 ;
      RECT  12.205 1.525 13.85 1.565 ;
      RECT  12.205 1.565 14.675 1.755 ;
      RECT  13.62 1.755 14.675 1.795 ;
      RECT  14.445 1.795 14.675 2.445 ;
      RECT  14.445 2.445 15.29 2.675 ;
      RECT  14.445 2.675 14.675 3.49 ;
      RECT  13.62 3.49 14.675 3.72 ;
      RECT  16.685 0.37 17.53 0.6 ;
      RECT  16.685 0.6 16.915 1.005 ;
      RECT  13.81 0.98 14.19 1.005 ;
      RECT  13.81 1.005 16.915 1.235 ;
      RECT  13.81 1.235 14.19 1.26 ;
      RECT  18.31 0.37 19.155 0.6 ;
      RECT  18.925 0.6 19.155 1.565 ;
      RECT  18.925 1.565 20.68 1.795 ;
      RECT  18.925 1.795 19.155 3.16 ;
      RECT  18.925 3.16 20.68 3.39 ;
      RECT  2.61 0.98 2.99 1.005 ;
      RECT  1.96 1.005 2.99 1.235 ;
      RECT  2.61 1.235 2.99 1.26 ;
      RECT  1.96 1.235 2.19 1.565 ;
      RECT  1.565 1.565 2.19 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 2.06 4.035 ;
      RECT  5.98 0.83 9.425 1.005 ;
      RECT  3.25 1.005 9.425 1.06 ;
      RECT  3.25 1.06 6.21 1.235 ;
      RECT  9.195 1.06 9.425 1.29 ;
      RECT  3.25 1.235 3.48 1.565 ;
      RECT  2.42 1.565 3.48 1.795 ;
      RECT  10.635 1.005 11.72 1.235 ;
      RECT  17.4 1.005 18.44 1.235 ;
      RECT  6.44 1.29 8.465 1.295 ;
      RECT  6.44 1.295 8.515 1.52 ;
      RECT  6.44 1.52 6.67 1.565 ;
      RECT  8.285 1.52 8.515 1.565 ;
      RECT  3.96 1.565 6.67 1.795 ;
      RECT  8.285 1.565 8.78 1.795 ;
      RECT  9.91 1.565 11.875 1.795 ;
      RECT  11.645 1.795 11.875 1.985 ;
      RECT  10.525 1.795 10.755 3.03 ;
      RECT  11.645 1.985 13.41 2.025 ;
      RECT  11.645 2.025 14.115 2.215 ;
      RECT  13.18 2.215 14.115 2.255 ;
      RECT  13.885 2.255 14.115 3.03 ;
      RECT  9.91 3.03 10.755 3.26 ;
      RECT  12.92 3.03 14.115 3.26 ;
      RECT  15.16 1.565 16.2 1.795 ;
      RECT  15.565 1.795 15.795 3.115 ;
      RECT  15.16 3.115 17.74 3.345 ;
      RECT  6.9 1.75 7.395 1.98 ;
      RECT  7.165 1.98 7.395 2.685 ;
      RECT  6.045 2.35 6.275 2.685 ;
      RECT  6.045 2.685 7.395 2.915 ;
      RECT  7.165 2.915 7.395 3.245 ;
      RECT  6.9 3.245 7.395 3.475 ;
      RECT  23.91 2.405 25.37 2.635 ;
      RECT  20.55 2.445 23.13 2.675 ;
      RECT  21.165 2.675 21.395 3.62 ;
      RECT  16.685 1.51 16.915 2.125 ;
      RECT  16.685 2.125 18.595 2.355 ;
      RECT  18.365 2.355 18.595 3.62 ;
      RECT  16.63 3.62 21.395 3.85 ;
      RECT  3.57 3.75 4.945 3.805 ;
      RECT  2.42 3.805 4.945 3.98 ;
      RECT  2.42 3.98 3.8 4.035 ;
      RECT  4.715 3.98 4.945 4.09 ;
      RECT  5.43 3.805 7.955 3.95 ;
      RECT  5.43 3.95 11.02 4.035 ;
      RECT  7.725 4.035 11.02 4.18 ;
      RECT  15.86 3.805 16.34 4.035 ;
      RECT  16.11 4.035 16.34 4.08 ;
      RECT  16.11 4.08 19.98 4.31 ;
      RECT  11.26 3.95 11.72 4.18 ;
      RECT  11.26 4.18 11.49 4.275 ;
      RECT  11.255 4.275 11.49 4.28 ;
      RECT  11.25 4.28 11.49 4.285 ;
      RECT  11.245 4.285 11.49 4.29 ;
      RECT  11.24 4.29 11.49 4.295 ;
      RECT  11.235 4.295 11.49 4.3 ;
      RECT  11.23 4.3 11.49 4.305 ;
      RECT  11.225 4.305 11.49 4.31 ;
      RECT  11.22 4.31 11.49 4.315 ;
      RECT  11.215 4.315 11.49 4.32 ;
      RECT  11.21 4.32 11.49 4.325 ;
      RECT  11.205 4.325 11.49 4.33 ;
      RECT  11.2 4.33 11.49 4.335 ;
      RECT  11.195 4.335 11.49 4.34 ;
      RECT  11.19 4.34 11.49 4.345 ;
      RECT  11.185 4.345 11.49 4.35 ;
      RECT  11.18 4.35 11.49 4.355 ;
      RECT  11.175 4.355 11.49 4.36 ;
      RECT  11.17 4.36 11.49 4.365 ;
      RECT  11.165 4.365 11.49 4.37 ;
      RECT  11.16 4.37 11.485 4.375 ;
      RECT  11.155 4.375 11.48 4.38 ;
      RECT  11.15 4.38 11.475 4.385 ;
      RECT  11.145 4.385 11.47 4.39 ;
      RECT  11.14 4.39 11.465 4.395 ;
      RECT  11.135 4.395 11.46 4.4 ;
      RECT  11.13 4.4 11.455 4.405 ;
      RECT  11.125 4.405 11.45 4.41 ;
      RECT  9.14 4.41 11.445 4.415 ;
      RECT  9.14 4.415 11.44 4.42 ;
      RECT  9.14 4.42 11.435 4.425 ;
      RECT  9.14 4.425 11.43 4.43 ;
      RECT  9.14 4.43 11.425 4.435 ;
      RECT  9.14 4.435 11.42 4.44 ;
      RECT  9.14 4.44 11.415 4.445 ;
      RECT  9.14 4.445 11.41 4.45 ;
      RECT  9.14 4.45 11.405 4.455 ;
      RECT  9.14 4.455 11.4 4.46 ;
      RECT  9.14 4.46 11.395 4.465 ;
      RECT  9.14 4.465 11.39 4.47 ;
      RECT  9.14 4.47 11.385 4.475 ;
      RECT  9.14 4.475 11.38 4.48 ;
      RECT  9.14 4.48 11.375 4.485 ;
      RECT  9.14 4.485 11.37 4.49 ;
      RECT  9.14 4.49 11.365 4.495 ;
      RECT  9.14 4.495 11.36 4.5 ;
      RECT  9.14 4.5 11.355 4.505 ;
      RECT  9.14 4.505 11.35 4.51 ;
      RECT  9.14 4.51 11.345 4.515 ;
      RECT  9.14 4.515 11.34 4.52 ;
      RECT  9.14 4.52 11.335 4.525 ;
      RECT  9.14 4.525 11.33 4.53 ;
      RECT  9.14 4.53 11.325 4.535 ;
      RECT  9.14 4.535 11.32 4.54 ;
      RECT  9.14 4.54 11.315 4.545 ;
      RECT  9.14 4.545 11.31 4.55 ;
      RECT  9.14 4.55 11.305 4.555 ;
      RECT  9.14 4.555 11.3 4.56 ;
      RECT  9.14 4.56 11.295 4.565 ;
      RECT  9.14 4.565 11.29 4.57 ;
      RECT  9.14 4.57 11.285 4.575 ;
      RECT  9.14 4.575 11.28 4.58 ;
      RECT  9.14 4.58 11.275 4.585 ;
      RECT  9.14 4.585 11.27 4.59 ;
      RECT  9.14 4.59 11.265 4.595 ;
      RECT  9.14 4.595 11.26 4.6 ;
      RECT  9.14 4.6 11.255 4.605 ;
      RECT  9.14 4.605 11.25 4.61 ;
      RECT  9.14 4.61 11.245 4.615 ;
      RECT  9.14 4.615 11.24 4.62 ;
      RECT  9.14 4.62 11.235 4.625 ;
      RECT  9.14 4.625 11.23 4.63 ;
      RECT  9.14 4.63 11.225 4.635 ;
      RECT  9.14 4.635 11.22 4.64 ;
      RECT  3.96 4.215 4.485 4.365 ;
      RECT  3.96 4.365 6.54 4.445 ;
      RECT  4.25 4.445 6.54 4.595 ;
      RECT  22.9 4.365 24.14 4.595 ;
      RECT  22.9 4.595 23.13 5.0 ;
      RECT  23.91 4.595 24.14 5.0 ;
      RECT  22.79 5.0 23.13 5.23 ;
      RECT  23.91 5.0 24.25 5.23 ;
      RECT  11.68 4.62 15.135 4.85 ;
      RECT  11.68 4.85 11.91 5.0 ;
      RECT  14.905 4.85 15.135 5.0 ;
      RECT  7.165 4.47 8.515 4.7 ;
      RECT  7.165 4.7 7.395 4.925 ;
      RECT  8.285 4.7 8.515 5.0 ;
      RECT  0.18 4.365 3.475 4.595 ;
      RECT  3.245 4.595 3.475 4.675 ;
      RECT  1.62 4.595 1.85 5.0 ;
      RECT  3.245 4.675 3.99 4.905 ;
      RECT  3.76 4.905 3.99 4.925 ;
      RECT  3.76 4.925 7.395 5.155 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  8.285 5.0 11.91 5.23 ;
      RECT  14.905 5.0 16.42 5.23 ;
      LAYER METAL2 ;
      RECT  2.61 0.98 14.19 1.26 ;
      LAYER VIA12 ;
      RECT  2.67 0.99 2.93 1.25 ;
      RECT  9.95 0.99 10.21 1.25 ;
      RECT  13.87 0.99 14.13 1.25 ;
  END
END MDN_FSDNRBQ_F_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNRBQ_1
#      Description : D-Flip Flop w/scan, neg-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNRBQ_1
  CLASS CORE ;
  FOREIGN MDN_FSDNRBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 1.565 2.94 2.695 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.485 1.565 19.98 1.795 ;
      RECT  19.485 1.795 19.715 3.245 ;
      RECT  19.485 3.245 19.98 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.98 2.125 16.38 2.355 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  14.445 5.08 14.675 5.46 ;
      RECT  12.88 5.46 14.675 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 10.64 5.74 ;
      RECT  5.43 5.085 5.77 5.46 ;
      RECT  5.04 5.46 6.16 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.565 ;
      RECT  15.12 -0.14 16.24 0.14 ;
      RECT  15.565 0.14 15.795 1.005 ;
      RECT  15.16 1.005 16.2 1.235 ;
      RECT  12.88 -0.14 14.0 0.14 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.52 ;
      RECT  3.805 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.6 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  10.425 0.37 13.05 0.6 ;
      RECT  10.425 0.6 10.655 0.75 ;
      RECT  5.98 0.37 9.635 0.6 ;
      RECT  9.405 0.6 9.635 0.75 ;
      RECT  5.98 0.6 6.21 0.83 ;
      RECT  9.405 0.75 10.655 0.98 ;
      RECT  4.715 0.83 6.21 1.06 ;
      RECT  4.715 1.06 4.945 1.29 ;
      RECT  19.43 0.37 19.77 0.6 ;
      RECT  19.43 0.6 19.66 0.795 ;
      RECT  18.31 0.37 18.65 0.6 ;
      RECT  18.42 0.6 18.65 0.795 ;
      RECT  18.42 0.795 19.66 1.025 ;
      RECT  6.44 0.83 8.78 1.06 ;
      RECT  8.44 1.06 8.78 1.12 ;
      RECT  6.44 1.06 6.67 1.29 ;
      RECT  5.485 1.29 6.67 1.52 ;
      RECT  5.485 1.52 5.715 1.565 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  3.245 1.565 5.715 1.795 ;
      RECT  10.885 0.83 13.96 1.06 ;
      RECT  13.62 1.06 13.96 1.12 ;
      RECT  10.885 1.06 11.115 1.235 ;
      RECT  8.995 1.235 11.115 1.24 ;
      RECT  8.99 1.24 11.115 1.245 ;
      RECT  8.985 1.245 11.115 1.25 ;
      RECT  8.98 1.25 11.115 1.255 ;
      RECT  8.975 1.255 11.115 1.26 ;
      RECT  8.97 1.26 11.115 1.265 ;
      RECT  8.965 1.265 11.115 1.27 ;
      RECT  8.96 1.27 11.115 1.275 ;
      RECT  8.955 1.275 11.115 1.28 ;
      RECT  8.95 1.28 11.115 1.285 ;
      RECT  8.945 1.285 11.115 1.29 ;
      RECT  8.94 1.29 11.115 1.295 ;
      RECT  8.935 1.295 11.115 1.3 ;
      RECT  8.93 1.3 11.115 1.305 ;
      RECT  8.925 1.305 11.115 1.31 ;
      RECT  8.92 1.31 11.115 1.315 ;
      RECT  8.915 1.315 11.115 1.32 ;
      RECT  8.91 1.32 11.115 1.325 ;
      RECT  8.905 1.325 11.115 1.33 ;
      RECT  8.9 1.33 11.115 1.335 ;
      RECT  8.895 1.335 11.115 1.34 ;
      RECT  8.89 1.34 11.115 1.345 ;
      RECT  8.885 1.345 11.115 1.35 ;
      RECT  6.9 1.29 8.265 1.295 ;
      RECT  6.9 1.295 8.27 1.3 ;
      RECT  6.9 1.3 8.275 1.305 ;
      RECT  6.9 1.305 8.28 1.31 ;
      RECT  6.9 1.31 8.285 1.315 ;
      RECT  6.9 1.315 8.29 1.32 ;
      RECT  6.9 1.32 8.295 1.325 ;
      RECT  6.9 1.325 8.3 1.33 ;
      RECT  6.9 1.33 8.305 1.335 ;
      RECT  6.9 1.335 8.31 1.34 ;
      RECT  6.9 1.34 8.315 1.345 ;
      RECT  6.9 1.345 8.32 1.35 ;
      RECT  6.9 1.35 11.115 1.465 ;
      RECT  6.9 1.465 9.09 1.47 ;
      RECT  6.9 1.47 9.085 1.475 ;
      RECT  6.9 1.475 9.08 1.48 ;
      RECT  6.9 1.48 9.075 1.485 ;
      RECT  6.9 1.485 9.07 1.49 ;
      RECT  6.9 1.49 9.065 1.495 ;
      RECT  6.9 1.495 9.06 1.5 ;
      RECT  6.9 1.5 9.055 1.505 ;
      RECT  6.9 1.505 9.05 1.51 ;
      RECT  6.9 1.51 9.045 1.515 ;
      RECT  6.9 1.515 9.04 1.52 ;
      RECT  8.16 1.52 9.035 1.525 ;
      RECT  8.165 1.525 9.03 1.53 ;
      RECT  8.17 1.53 9.025 1.535 ;
      RECT  8.175 1.535 9.02 1.54 ;
      RECT  8.18 1.54 9.015 1.545 ;
      RECT  8.185 1.545 9.01 1.55 ;
      RECT  8.19 1.55 9.005 1.555 ;
      RECT  8.195 1.555 9.0 1.56 ;
      RECT  8.2 1.56 8.995 1.565 ;
      RECT  8.205 1.565 8.99 1.57 ;
      RECT  8.21 1.57 8.985 1.575 ;
      RECT  8.215 1.575 8.98 1.58 ;
      RECT  16.685 1.005 18.035 1.235 ;
      RECT  17.805 1.235 18.035 1.255 ;
      RECT  16.685 1.235 16.915 1.565 ;
      RECT  17.805 1.255 18.385 1.485 ;
      RECT  18.155 1.485 18.385 1.85 ;
      RECT  11.38 1.29 13.465 1.295 ;
      RECT  11.38 1.295 13.47 1.3 ;
      RECT  11.38 1.3 13.475 1.305 ;
      RECT  11.38 1.305 13.48 1.31 ;
      RECT  11.38 1.31 13.485 1.315 ;
      RECT  11.38 1.315 13.49 1.32 ;
      RECT  11.38 1.32 13.495 1.325 ;
      RECT  11.38 1.325 13.5 1.33 ;
      RECT  11.38 1.33 13.505 1.335 ;
      RECT  11.38 1.335 13.51 1.34 ;
      RECT  11.38 1.34 13.515 1.345 ;
      RECT  11.38 1.345 13.52 1.35 ;
      RECT  11.38 1.35 13.525 1.355 ;
      RECT  11.38 1.355 13.53 1.36 ;
      RECT  11.38 1.36 13.535 1.365 ;
      RECT  11.38 1.365 13.54 1.37 ;
      RECT  11.38 1.37 13.545 1.375 ;
      RECT  11.38 1.375 13.55 1.38 ;
      RECT  11.38 1.38 13.555 1.385 ;
      RECT  11.38 1.385 13.56 1.39 ;
      RECT  11.38 1.39 13.565 1.395 ;
      RECT  11.38 1.395 13.57 1.4 ;
      RECT  11.38 1.4 13.575 1.405 ;
      RECT  11.38 1.405 13.58 1.41 ;
      RECT  11.38 1.41 13.585 1.415 ;
      RECT  11.38 1.415 13.59 1.42 ;
      RECT  11.38 1.42 13.595 1.425 ;
      RECT  11.38 1.425 13.6 1.43 ;
      RECT  11.38 1.43 13.605 1.435 ;
      RECT  11.38 1.435 13.61 1.44 ;
      RECT  11.38 1.44 13.615 1.445 ;
      RECT  11.38 1.445 13.62 1.45 ;
      RECT  11.38 1.45 13.625 1.455 ;
      RECT  11.38 1.455 13.63 1.46 ;
      RECT  11.38 1.46 13.635 1.465 ;
      RECT  11.38 1.465 13.64 1.47 ;
      RECT  11.38 1.47 13.645 1.475 ;
      RECT  11.38 1.475 13.65 1.48 ;
      RECT  11.38 1.48 13.655 1.485 ;
      RECT  11.38 1.485 13.66 1.49 ;
      RECT  11.38 1.49 13.665 1.495 ;
      RECT  11.38 1.495 13.67 1.5 ;
      RECT  11.38 1.5 13.675 1.505 ;
      RECT  11.38 1.505 13.68 1.51 ;
      RECT  11.38 1.51 13.685 1.515 ;
      RECT  11.38 1.515 13.69 1.52 ;
      RECT  13.36 1.52 13.695 1.525 ;
      RECT  13.365 1.525 13.7 1.53 ;
      RECT  13.37 1.53 13.705 1.535 ;
      RECT  13.375 1.535 13.71 1.54 ;
      RECT  13.38 1.54 13.715 1.545 ;
      RECT  13.385 1.545 13.72 1.55 ;
      RECT  13.39 1.55 13.725 1.555 ;
      RECT  13.395 1.555 13.73 1.56 ;
      RECT  13.4 1.56 13.735 1.565 ;
      RECT  13.405 1.565 16.915 1.57 ;
      RECT  13.41 1.57 16.915 1.575 ;
      RECT  13.415 1.575 16.915 1.58 ;
      RECT  13.42 1.58 16.915 1.585 ;
      RECT  13.425 1.585 16.915 1.59 ;
      RECT  13.43 1.59 16.915 1.595 ;
      RECT  13.435 1.595 16.915 1.6 ;
      RECT  13.44 1.6 16.915 1.605 ;
      RECT  13.445 1.605 16.915 1.61 ;
      RECT  13.45 1.61 16.915 1.615 ;
      RECT  13.455 1.615 16.915 1.62 ;
      RECT  13.46 1.62 16.915 1.625 ;
      RECT  13.465 1.625 16.915 1.63 ;
      RECT  13.47 1.63 16.915 1.635 ;
      RECT  13.475 1.635 16.915 1.64 ;
      RECT  13.48 1.64 16.915 1.645 ;
      RECT  13.485 1.645 16.915 1.65 ;
      RECT  13.49 1.65 16.915 1.655 ;
      RECT  13.495 1.655 16.915 1.66 ;
      RECT  13.5 1.66 16.915 1.665 ;
      RECT  13.505 1.665 16.915 1.67 ;
      RECT  13.51 1.67 16.915 1.675 ;
      RECT  13.515 1.675 16.915 1.68 ;
      RECT  13.52 1.68 16.915 1.685 ;
      RECT  13.525 1.685 16.915 1.69 ;
      RECT  13.53 1.69 16.915 1.695 ;
      RECT  13.535 1.695 16.915 1.7 ;
      RECT  13.54 1.7 16.915 1.705 ;
      RECT  13.545 1.705 16.915 1.71 ;
      RECT  13.55 1.71 16.915 1.715 ;
      RECT  13.555 1.715 16.915 1.72 ;
      RECT  13.56 1.72 16.915 1.725 ;
      RECT  13.565 1.725 16.915 1.73 ;
      RECT  13.57 1.73 16.915 1.735 ;
      RECT  13.575 1.735 16.915 1.74 ;
      RECT  13.58 1.74 16.915 1.745 ;
      RECT  13.585 1.745 16.915 1.75 ;
      RECT  13.59 1.75 16.915 1.755 ;
      RECT  13.595 1.755 16.915 1.76 ;
      RECT  13.6 1.76 16.915 1.765 ;
      RECT  13.605 1.765 16.915 1.77 ;
      RECT  13.61 1.77 16.915 1.775 ;
      RECT  13.615 1.775 16.915 1.78 ;
      RECT  13.62 1.78 16.915 1.785 ;
      RECT  13.625 1.785 16.915 1.79 ;
      RECT  13.63 1.79 16.915 1.795 ;
      RECT  7.62 1.75 7.96 1.82 ;
      RECT  7.62 1.82 8.91 2.05 ;
      RECT  8.68 2.05 8.91 2.66 ;
      RECT  8.68 2.66 9.15 2.835 ;
      RECT  7.725 2.835 9.15 2.94 ;
      RECT  7.725 2.94 8.91 3.065 ;
      RECT  7.725 3.065 7.955 3.315 ;
      RECT  17.4 1.715 17.74 1.945 ;
      RECT  17.51 1.945 17.74 2.125 ;
      RECT  17.51 2.125 18.595 2.355 ;
      RECT  18.365 2.355 18.595 3.245 ;
      RECT  15.86 3.245 18.595 3.475 ;
      RECT  6.2 1.75 6.835 1.98 ;
      RECT  6.605 1.98 6.835 2.365 ;
      RECT  6.605 2.365 8.45 2.595 ;
      RECT  6.605 2.595 6.835 3.245 ;
      RECT  6.2 3.245 6.835 3.475 ;
      RECT  9.14 1.75 10.195 1.98 ;
      RECT  9.965 1.98 10.195 3.755 ;
      RECT  8.645 3.755 10.195 3.985 ;
      RECT  8.645 3.985 8.875 4.02 ;
      RECT  7.725 4.02 8.875 4.25 ;
      RECT  7.725 4.25 7.955 4.925 ;
      RECT  4.925 4.625 6.275 4.855 ;
      RECT  6.045 4.855 6.275 4.925 ;
      RECT  4.925 4.855 5.155 5.0 ;
      RECT  6.045 4.925 7.955 5.155 ;
      RECT  3.75 5.0 5.155 5.23 ;
      RECT  12.15 1.75 12.49 1.98 ;
      RECT  12.205 1.98 12.435 3.315 ;
      RECT  12.765 1.75 13.26 1.98 ;
      RECT  12.765 1.98 12.995 2.685 ;
      RECT  12.665 2.685 14.115 2.915 ;
      RECT  13.885 2.35 14.115 2.685 ;
      RECT  12.665 2.915 12.895 3.545 ;
      RECT  10.68 1.75 11.315 1.98 ;
      RECT  11.085 1.98 11.315 3.545 ;
      RECT  10.68 3.545 12.895 3.775 ;
      RECT  10.47 2.34 10.81 2.66 ;
      RECT  10.43 2.66 10.81 2.94 ;
      RECT  6.045 2.35 6.275 2.685 ;
      RECT  5.485 2.685 6.275 2.915 ;
      RECT  5.485 2.915 5.715 3.245 ;
      RECT  4.66 3.245 5.715 3.475 ;
      RECT  9.405 2.35 9.635 3.295 ;
      RECT  8.185 3.295 9.635 3.525 ;
      RECT  8.185 3.525 8.415 3.56 ;
      RECT  7.165 3.56 8.415 3.705 ;
      RECT  3.805 3.705 8.415 3.79 ;
      RECT  3.805 3.79 7.395 3.935 ;
      RECT  3.805 3.935 4.035 4.08 ;
      RECT  2.685 4.08 4.035 4.31 ;
      RECT  2.685 4.31 2.915 4.925 ;
      RECT  1.51 4.925 2.915 5.155 ;
      RECT  1.51 5.155 1.85 5.23 ;
      RECT  1.72 3.145 2.76 3.375 ;
      RECT  3.245 3.245 4.3 3.475 ;
      RECT  3.245 3.475 3.475 3.605 ;
      RECT  2.125 3.605 3.475 3.835 ;
      RECT  2.125 3.835 2.355 4.365 ;
      RECT  0.18 4.365 2.355 4.595 ;
      RECT  13.125 3.245 15.5 3.475 ;
      RECT  13.125 3.475 13.355 4.005 ;
      RECT  12.205 4.005 13.355 4.215 ;
      RECT  9.105 4.215 13.355 4.235 ;
      RECT  9.105 4.235 12.435 4.445 ;
      RECT  9.105 4.445 9.335 4.48 ;
      RECT  8.44 4.48 9.335 4.71 ;
      RECT  13.585 3.805 18.44 4.035 ;
      RECT  13.585 4.035 13.815 4.465 ;
      RECT  12.92 4.465 13.815 4.695 ;
      RECT  4.365 4.165 7.24 4.395 ;
      RECT  4.365 4.395 4.595 4.54 ;
      RECT  3.245 4.54 4.595 4.77 ;
      RECT  3.245 4.77 3.475 5.21 ;
      RECT  14.045 4.365 17.41 4.595 ;
      RECT  14.045 4.595 14.275 4.825 ;
      RECT  17.18 4.595 17.41 5.0 ;
      RECT  14.04 4.825 14.275 4.83 ;
      RECT  14.035 4.83 14.275 4.835 ;
      RECT  14.03 4.835 14.275 4.84 ;
      RECT  14.025 4.84 14.275 4.845 ;
      RECT  14.02 4.845 14.275 4.85 ;
      RECT  14.015 4.85 14.275 4.855 ;
      RECT  14.01 4.855 14.275 4.86 ;
      RECT  14.005 4.86 14.275 4.865 ;
      RECT  14.0 4.865 14.275 4.87 ;
      RECT  13.995 4.87 14.275 4.875 ;
      RECT  13.99 4.875 14.275 4.88 ;
      RECT  13.985 4.88 14.275 4.885 ;
      RECT  13.98 4.885 14.275 4.89 ;
      RECT  13.975 4.89 14.275 4.895 ;
      RECT  13.97 4.895 14.275 4.9 ;
      RECT  13.965 4.9 14.275 4.905 ;
      RECT  13.96 4.905 14.275 4.91 ;
      RECT  13.955 4.91 14.275 4.915 ;
      RECT  13.95 4.915 14.275 4.92 ;
      RECT  13.945 4.92 14.27 4.925 ;
      RECT  12.15 4.925 14.265 4.93 ;
      RECT  12.15 4.93 14.26 4.935 ;
      RECT  12.15 4.935 14.255 4.94 ;
      RECT  12.15 4.94 14.25 4.945 ;
      RECT  12.15 4.945 14.245 4.95 ;
      RECT  12.15 4.95 14.24 4.955 ;
      RECT  12.15 4.955 14.235 4.96 ;
      RECT  12.15 4.96 14.23 4.965 ;
      RECT  12.15 4.965 14.225 4.97 ;
      RECT  12.15 4.97 14.22 4.975 ;
      RECT  12.15 4.975 14.215 4.98 ;
      RECT  12.15 4.98 14.21 4.985 ;
      RECT  12.15 4.985 14.205 4.99 ;
      RECT  12.15 4.99 14.2 4.995 ;
      RECT  12.15 4.995 14.195 5.0 ;
      RECT  12.15 5.0 14.19 5.005 ;
      RECT  17.18 5.0 17.53 5.23 ;
      RECT  12.15 5.005 14.185 5.01 ;
      RECT  12.15 5.01 14.18 5.015 ;
      RECT  12.15 5.015 14.175 5.02 ;
      RECT  12.15 5.02 14.17 5.025 ;
      RECT  12.15 5.025 14.165 5.03 ;
      RECT  12.15 5.03 14.16 5.035 ;
      RECT  12.15 5.035 14.155 5.04 ;
      RECT  12.15 5.04 14.15 5.045 ;
      RECT  12.15 5.045 14.145 5.05 ;
      RECT  12.15 5.05 14.14 5.055 ;
      RECT  12.15 5.055 14.135 5.06 ;
      RECT  12.15 5.06 14.13 5.065 ;
      RECT  12.15 5.065 14.125 5.07 ;
      RECT  12.15 5.07 14.12 5.075 ;
      RECT  12.15 5.075 14.115 5.08 ;
      RECT  12.15 5.08 14.11 5.085 ;
      RECT  12.15 5.085 14.105 5.09 ;
      RECT  12.15 5.09 14.1 5.095 ;
      RECT  12.15 5.095 14.095 5.1 ;
      RECT  12.15 5.1 14.09 5.105 ;
      RECT  12.15 5.105 14.085 5.11 ;
      RECT  12.15 5.11 14.08 5.115 ;
      RECT  12.15 5.115 14.075 5.12 ;
      RECT  12.15 5.12 14.07 5.125 ;
      RECT  12.15 5.125 14.065 5.13 ;
      RECT  12.15 5.13 14.06 5.135 ;
      RECT  12.15 5.135 14.055 5.14 ;
      RECT  12.15 5.14 14.05 5.145 ;
      RECT  12.15 5.145 14.045 5.15 ;
      RECT  12.15 5.15 14.04 5.155 ;
      RECT  9.71 4.675 10.755 4.68 ;
      RECT  9.705 4.68 10.755 4.685 ;
      RECT  9.7 4.685 10.755 4.69 ;
      RECT  9.695 4.69 10.755 4.695 ;
      RECT  9.69 4.695 10.755 4.7 ;
      RECT  9.685 4.7 10.755 4.705 ;
      RECT  9.68 4.705 10.755 4.71 ;
      RECT  9.675 4.71 10.755 4.715 ;
      RECT  9.67 4.715 10.755 4.72 ;
      RECT  9.665 4.72 10.755 4.725 ;
      RECT  9.66 4.725 10.755 4.73 ;
      RECT  9.655 4.73 10.755 4.735 ;
      RECT  9.65 4.735 10.755 4.74 ;
      RECT  9.645 4.74 10.755 4.745 ;
      RECT  9.64 4.745 10.755 4.75 ;
      RECT  9.635 4.75 10.755 4.755 ;
      RECT  9.63 4.755 10.755 4.76 ;
      RECT  9.625 4.76 10.755 4.765 ;
      RECT  9.62 4.765 10.755 4.77 ;
      RECT  9.615 4.77 10.755 4.775 ;
      RECT  9.61 4.775 10.755 4.78 ;
      RECT  9.605 4.78 10.755 4.785 ;
      RECT  9.6 4.785 10.755 4.79 ;
      RECT  9.595 4.79 10.755 4.795 ;
      RECT  9.59 4.795 10.755 4.8 ;
      RECT  9.585 4.8 10.755 4.805 ;
      RECT  9.58 4.805 10.755 4.81 ;
      RECT  9.575 4.81 10.755 4.815 ;
      RECT  9.57 4.815 10.755 4.82 ;
      RECT  9.565 4.82 10.755 4.825 ;
      RECT  9.56 4.825 10.755 4.83 ;
      RECT  9.555 4.83 10.755 4.835 ;
      RECT  9.55 4.835 10.755 4.84 ;
      RECT  9.545 4.84 10.755 4.845 ;
      RECT  9.54 4.845 10.755 4.85 ;
      RECT  9.535 4.85 10.755 4.855 ;
      RECT  9.53 4.855 10.755 4.86 ;
      RECT  9.525 4.86 10.755 4.865 ;
      RECT  9.52 4.865 10.755 4.87 ;
      RECT  9.515 4.87 10.755 4.875 ;
      RECT  9.51 4.875 10.755 4.88 ;
      RECT  9.505 4.88 10.755 4.885 ;
      RECT  9.5 4.885 10.755 4.89 ;
      RECT  9.495 4.89 10.755 4.895 ;
      RECT  9.49 4.895 10.755 4.9 ;
      RECT  9.485 4.9 10.755 4.905 ;
      RECT  9.48 4.905 9.805 4.91 ;
      RECT  10.525 4.905 10.755 5.0 ;
      RECT  9.475 4.91 9.8 4.915 ;
      RECT  9.47 4.915 9.795 4.92 ;
      RECT  9.465 4.92 9.79 4.925 ;
      RECT  9.46 4.925 9.785 4.93 ;
      RECT  9.455 4.93 9.78 4.935 ;
      RECT  9.45 4.935 9.775 4.94 ;
      RECT  9.445 4.94 9.77 4.945 ;
      RECT  9.44 4.945 9.765 4.95 ;
      RECT  9.435 4.95 9.76 4.955 ;
      RECT  9.43 4.955 9.755 4.96 ;
      RECT  9.425 4.96 9.75 4.965 ;
      RECT  9.42 4.965 9.745 4.97 ;
      RECT  9.415 4.97 9.74 4.975 ;
      RECT  9.41 4.975 9.735 4.98 ;
      RECT  9.405 4.98 9.73 4.985 ;
      RECT  9.4 4.985 9.725 4.99 ;
      RECT  9.395 4.99 9.72 4.995 ;
      RECT  9.39 4.995 9.715 5.0 ;
      RECT  8.23 5.0 9.71 5.005 ;
      RECT  10.525 5.0 11.92 5.23 ;
      RECT  8.23 5.005 9.705 5.01 ;
      RECT  8.23 5.01 9.7 5.015 ;
      RECT  8.23 5.015 9.695 5.02 ;
      RECT  8.23 5.02 9.69 5.025 ;
      RECT  8.23 5.025 9.685 5.03 ;
      RECT  8.23 5.03 9.68 5.035 ;
      RECT  8.23 5.035 9.675 5.04 ;
      RECT  8.23 5.04 9.67 5.045 ;
      RECT  8.23 5.045 9.665 5.05 ;
      RECT  8.23 5.05 9.66 5.055 ;
      RECT  8.23 5.055 9.655 5.06 ;
      RECT  8.23 5.06 9.65 5.065 ;
      RECT  8.23 5.065 9.645 5.07 ;
      RECT  8.23 5.07 9.64 5.075 ;
      RECT  8.23 5.075 9.635 5.08 ;
      RECT  8.23 5.08 9.63 5.085 ;
      RECT  8.23 5.085 9.625 5.09 ;
      RECT  8.23 5.09 9.62 5.095 ;
      RECT  8.23 5.095 9.615 5.1 ;
      RECT  8.23 5.1 9.61 5.105 ;
      RECT  8.23 5.105 9.605 5.11 ;
      RECT  8.23 5.11 9.6 5.115 ;
      RECT  8.23 5.115 9.595 5.12 ;
      RECT  8.23 5.12 9.59 5.125 ;
      RECT  8.23 5.125 9.585 5.13 ;
      RECT  8.23 5.13 9.58 5.135 ;
      RECT  8.23 5.135 9.575 5.14 ;
      RECT  8.23 5.14 9.57 5.145 ;
      RECT  8.23 5.145 9.565 5.15 ;
      RECT  8.23 5.15 9.56 5.155 ;
      RECT  8.23 5.155 9.555 5.16 ;
      RECT  8.23 5.16 9.55 5.165 ;
      RECT  8.23 5.165 9.545 5.17 ;
      RECT  8.23 5.17 9.54 5.175 ;
      RECT  8.23 5.175 9.535 5.18 ;
      RECT  8.23 5.18 9.53 5.185 ;
      RECT  8.23 5.185 9.525 5.19 ;
      RECT  8.23 5.19 9.52 5.195 ;
      RECT  8.23 5.195 9.515 5.2 ;
      RECT  8.23 5.2 9.51 5.205 ;
      RECT  8.23 5.205 9.505 5.21 ;
      RECT  8.23 5.21 9.5 5.215 ;
      RECT  8.23 5.215 9.495 5.22 ;
      RECT  8.23 5.22 9.49 5.225 ;
      RECT  8.23 5.225 9.485 5.23 ;
      LAYER METAL2 ;
      RECT  8.77 2.66 10.81 2.94 ;
      LAYER VIA12 ;
      RECT  8.83 2.67 9.09 2.93 ;
      RECT  10.49 2.67 10.75 2.93 ;
  END
END MDN_FSDNRBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNRBQ_2
#      Description : D-Flip Flop w/scan, neg-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNRBQ_2
  CLASS CORE ;
  FOREIGN MDN_FSDNRBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 1.565 2.94 2.69 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.64 1.565 20.68 1.795 ;
      RECT  20.045 1.795 20.275 3.245 ;
      RECT  19.64 3.245 20.685 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.98 2.125 16.38 2.355 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.405 2.35 9.635 3.26 ;
      RECT  8.2 3.26 9.635 3.49 ;
      RECT  8.2 3.49 8.43 3.545 ;
      RECT  7.165 3.5 7.47 3.545 ;
      RECT  7.165 3.545 8.43 3.755 ;
      RECT  3.73 3.755 8.43 3.775 ;
      RECT  3.73 3.775 7.47 3.985 ;
      RECT  3.73 3.985 4.035 4.08 ;
      RECT  2.685 4.08 4.035 4.31 ;
      RECT  2.685 4.31 2.99 4.365 ;
      RECT  1.51 4.365 2.99 4.595 ;
      RECT  1.51 4.595 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  14.445 5.08 14.675 5.46 ;
      RECT  12.88 5.46 14.675 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 10.64 5.74 ;
      RECT  5.43 5.135 5.77 5.46 ;
      RECT  5.04 5.46 6.16 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 22.57 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  15.12 -0.14 16.24 0.14 ;
      RECT  15.565 0.14 15.795 1.005 ;
      RECT  15.16 1.005 16.2 1.235 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.6 ;
      RECT  3.805 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.6 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  20.31 -0.13 20.57 0.13 ;
      RECT  20.87 -0.13 21.13 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  10.425 0.37 13.05 0.6 ;
      RECT  10.425 0.6 10.655 0.83 ;
      RECT  5.98 0.37 9.635 0.6 ;
      RECT  5.98 0.6 6.21 0.83 ;
      RECT  9.405 0.6 9.635 0.83 ;
      RECT  4.715 0.83 6.21 1.06 ;
      RECT  9.405 0.83 10.655 1.06 ;
      RECT  4.715 1.06 4.945 1.29 ;
      RECT  19.43 0.37 20.89 0.6 ;
      RECT  10.885 0.83 13.955 0.89 ;
      RECT  10.885 0.89 13.96 1.06 ;
      RECT  13.62 1.06 13.96 1.12 ;
      RECT  10.885 1.06 11.115 1.29 ;
      RECT  8.94 1.29 11.115 1.295 ;
      RECT  8.935 1.295 11.115 1.3 ;
      RECT  8.93 1.3 11.115 1.305 ;
      RECT  8.925 1.305 11.115 1.31 ;
      RECT  8.92 1.31 11.115 1.315 ;
      RECT  8.915 1.315 11.115 1.32 ;
      RECT  8.91 1.32 11.115 1.325 ;
      RECT  8.905 1.325 11.115 1.33 ;
      RECT  8.9 1.33 11.115 1.335 ;
      RECT  8.895 1.335 11.115 1.34 ;
      RECT  8.89 1.34 11.115 1.345 ;
      RECT  8.885 1.345 11.115 1.35 ;
      RECT  6.9 1.29 8.22 1.295 ;
      RECT  6.9 1.295 8.225 1.3 ;
      RECT  6.9 1.3 8.23 1.305 ;
      RECT  6.9 1.305 8.235 1.31 ;
      RECT  6.9 1.31 8.24 1.315 ;
      RECT  6.9 1.315 8.245 1.32 ;
      RECT  6.9 1.32 8.25 1.325 ;
      RECT  6.9 1.325 8.255 1.33 ;
      RECT  6.9 1.33 8.26 1.335 ;
      RECT  6.9 1.335 8.265 1.34 ;
      RECT  6.9 1.34 8.27 1.345 ;
      RECT  6.9 1.345 8.275 1.35 ;
      RECT  6.9 1.35 11.115 1.52 ;
      RECT  8.115 1.52 9.035 1.525 ;
      RECT  8.12 1.525 9.03 1.53 ;
      RECT  8.125 1.53 9.025 1.535 ;
      RECT  8.13 1.535 9.02 1.54 ;
      RECT  8.135 1.54 9.015 1.545 ;
      RECT  8.14 1.545 9.01 1.55 ;
      RECT  8.145 1.55 9.005 1.555 ;
      RECT  8.15 1.555 9.0 1.56 ;
      RECT  8.155 1.56 8.995 1.565 ;
      RECT  8.16 1.565 8.99 1.57 ;
      RECT  8.165 1.57 8.985 1.575 ;
      RECT  8.17 1.575 8.98 1.58 ;
      RECT  6.44 0.83 8.78 1.06 ;
      RECT  8.44 1.06 8.78 1.12 ;
      RECT  6.44 1.06 6.67 1.29 ;
      RECT  5.485 1.29 6.67 1.52 ;
      RECT  5.485 1.52 5.715 1.565 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  3.245 1.565 5.715 1.795 ;
      RECT  16.685 1.005 18.445 1.235 ;
      RECT  16.685 1.235 16.915 1.565 ;
      RECT  11.38 1.29 13.465 1.295 ;
      RECT  11.38 1.295 13.47 1.3 ;
      RECT  11.38 1.3 13.475 1.305 ;
      RECT  11.38 1.305 13.48 1.31 ;
      RECT  11.38 1.31 13.485 1.315 ;
      RECT  11.38 1.315 13.49 1.32 ;
      RECT  11.38 1.32 13.495 1.325 ;
      RECT  11.38 1.325 13.5 1.33 ;
      RECT  11.38 1.33 13.505 1.335 ;
      RECT  11.38 1.335 13.51 1.34 ;
      RECT  11.38 1.34 13.515 1.345 ;
      RECT  11.38 1.345 13.52 1.35 ;
      RECT  11.38 1.35 13.525 1.355 ;
      RECT  11.38 1.355 13.53 1.36 ;
      RECT  11.38 1.36 13.535 1.365 ;
      RECT  11.38 1.365 13.54 1.37 ;
      RECT  11.38 1.37 13.545 1.375 ;
      RECT  11.38 1.375 13.55 1.38 ;
      RECT  11.38 1.38 13.555 1.385 ;
      RECT  11.38 1.385 13.56 1.39 ;
      RECT  11.38 1.39 13.565 1.395 ;
      RECT  11.38 1.395 13.57 1.4 ;
      RECT  11.38 1.4 13.575 1.405 ;
      RECT  11.38 1.405 13.58 1.41 ;
      RECT  11.38 1.41 13.585 1.415 ;
      RECT  11.38 1.415 13.59 1.42 ;
      RECT  11.38 1.42 13.595 1.425 ;
      RECT  11.38 1.425 13.6 1.43 ;
      RECT  11.38 1.43 13.605 1.435 ;
      RECT  11.38 1.435 13.61 1.44 ;
      RECT  11.38 1.44 13.615 1.445 ;
      RECT  11.38 1.445 13.62 1.45 ;
      RECT  11.38 1.45 13.625 1.455 ;
      RECT  11.38 1.455 13.63 1.46 ;
      RECT  11.38 1.46 13.635 1.465 ;
      RECT  11.38 1.465 13.64 1.47 ;
      RECT  11.38 1.47 13.645 1.475 ;
      RECT  11.38 1.475 13.65 1.48 ;
      RECT  11.38 1.48 13.655 1.485 ;
      RECT  11.38 1.485 13.66 1.49 ;
      RECT  11.38 1.49 13.665 1.495 ;
      RECT  11.38 1.495 13.67 1.5 ;
      RECT  11.38 1.5 13.675 1.505 ;
      RECT  11.38 1.505 13.68 1.51 ;
      RECT  11.38 1.51 13.685 1.515 ;
      RECT  11.38 1.515 13.69 1.52 ;
      RECT  13.36 1.52 13.695 1.525 ;
      RECT  13.365 1.525 13.7 1.53 ;
      RECT  13.37 1.53 13.705 1.535 ;
      RECT  13.375 1.535 13.71 1.54 ;
      RECT  13.38 1.54 13.715 1.545 ;
      RECT  13.385 1.545 13.72 1.55 ;
      RECT  13.39 1.55 13.725 1.555 ;
      RECT  13.395 1.555 13.73 1.56 ;
      RECT  13.4 1.56 13.735 1.565 ;
      RECT  13.405 1.565 16.92 1.57 ;
      RECT  13.41 1.57 16.92 1.575 ;
      RECT  13.415 1.575 16.92 1.58 ;
      RECT  13.42 1.58 16.92 1.585 ;
      RECT  13.425 1.585 16.92 1.59 ;
      RECT  13.43 1.59 16.92 1.595 ;
      RECT  13.435 1.595 16.92 1.6 ;
      RECT  13.44 1.6 16.92 1.605 ;
      RECT  13.445 1.605 16.92 1.61 ;
      RECT  13.45 1.61 16.92 1.615 ;
      RECT  13.455 1.615 16.92 1.62 ;
      RECT  13.46 1.62 16.92 1.625 ;
      RECT  13.465 1.625 16.92 1.63 ;
      RECT  13.47 1.63 16.92 1.635 ;
      RECT  13.475 1.635 16.92 1.64 ;
      RECT  13.48 1.64 16.92 1.645 ;
      RECT  13.485 1.645 16.92 1.65 ;
      RECT  13.49 1.65 16.92 1.655 ;
      RECT  13.495 1.655 16.92 1.66 ;
      RECT  13.5 1.66 16.92 1.665 ;
      RECT  13.505 1.665 16.92 1.67 ;
      RECT  13.51 1.67 16.92 1.675 ;
      RECT  13.515 1.675 16.92 1.68 ;
      RECT  13.52 1.68 16.92 1.685 ;
      RECT  13.525 1.685 16.92 1.69 ;
      RECT  13.53 1.69 16.92 1.695 ;
      RECT  13.535 1.695 16.92 1.7 ;
      RECT  13.54 1.7 16.92 1.705 ;
      RECT  13.545 1.705 16.92 1.71 ;
      RECT  13.55 1.71 16.92 1.715 ;
      RECT  13.555 1.715 16.92 1.72 ;
      RECT  13.56 1.72 16.92 1.725 ;
      RECT  13.565 1.725 16.92 1.73 ;
      RECT  13.57 1.73 16.92 1.735 ;
      RECT  13.575 1.735 16.92 1.74 ;
      RECT  13.58 1.74 16.92 1.745 ;
      RECT  13.585 1.745 16.92 1.75 ;
      RECT  13.59 1.75 16.92 1.755 ;
      RECT  13.595 1.755 16.92 1.76 ;
      RECT  13.6 1.76 16.92 1.765 ;
      RECT  13.605 1.765 16.92 1.77 ;
      RECT  13.61 1.77 16.92 1.775 ;
      RECT  13.615 1.775 16.92 1.78 ;
      RECT  13.62 1.78 16.92 1.785 ;
      RECT  13.625 1.785 16.92 1.79 ;
      RECT  13.63 1.79 16.92 1.795 ;
      RECT  17.4 1.565 18.595 1.795 ;
      RECT  18.365 1.795 18.595 2.685 ;
      RECT  18.365 2.685 19.715 2.915 ;
      RECT  19.485 2.355 19.715 2.685 ;
      RECT  18.365 2.915 18.595 3.245 ;
      RECT  15.86 3.245 18.595 3.475 ;
      RECT  7.63 1.75 7.97 1.82 ;
      RECT  7.63 1.82 8.865 2.05 ;
      RECT  8.635 2.05 8.865 2.66 ;
      RECT  8.635 2.66 9.15 2.8 ;
      RECT  7.725 2.8 9.15 2.94 ;
      RECT  7.725 2.94 8.865 3.03 ;
      RECT  7.725 3.03 7.955 3.315 ;
      RECT  6.2 1.75 6.835 1.98 ;
      RECT  6.605 1.98 6.835 2.34 ;
      RECT  6.605 2.34 8.405 2.57 ;
      RECT  6.605 2.57 6.835 3.245 ;
      RECT  6.2 3.245 6.835 3.475 ;
      RECT  9.14 1.75 10.195 1.98 ;
      RECT  9.965 1.98 10.195 3.72 ;
      RECT  8.66 3.72 10.195 3.95 ;
      RECT  8.66 3.95 8.89 4.005 ;
      RECT  7.725 4.005 8.89 4.235 ;
      RECT  7.725 4.235 7.955 4.925 ;
      RECT  4.925 4.675 6.275 4.905 ;
      RECT  6.045 4.905 6.275 4.925 ;
      RECT  4.925 4.905 5.155 5.0 ;
      RECT  6.045 4.925 7.955 5.155 ;
      RECT  3.75 5.0 5.155 5.23 ;
      RECT  12.15 1.75 12.49 1.98 ;
      RECT  12.15 1.98 12.38 2.975 ;
      RECT  12.15 2.975 12.435 3.315 ;
      RECT  12.765 1.75 13.26 1.98 ;
      RECT  12.765 1.98 12.995 2.685 ;
      RECT  12.665 2.685 14.115 2.915 ;
      RECT  13.885 2.39 14.115 2.685 ;
      RECT  12.665 2.915 12.895 3.545 ;
      RECT  10.68 1.75 11.315 1.98 ;
      RECT  11.085 1.98 11.315 3.545 ;
      RECT  10.68 3.545 12.895 3.775 ;
      RECT  5.485 2.41 6.33 2.64 ;
      RECT  5.485 2.64 5.715 3.245 ;
      RECT  4.66 3.245 5.715 3.475 ;
      RECT  10.47 2.28 10.81 2.66 ;
      RECT  10.45 2.66 10.83 2.94 ;
      RECT  1.72 3.16 2.76 3.39 ;
      RECT  3.245 3.245 4.3 3.475 ;
      RECT  3.245 3.475 3.475 3.62 ;
      RECT  2.125 3.62 3.475 3.805 ;
      RECT  0.18 3.805 3.475 3.85 ;
      RECT  0.18 3.85 2.355 4.035 ;
      RECT  13.125 3.245 15.5 3.475 ;
      RECT  13.125 3.475 13.355 4.005 ;
      RECT  12.205 4.005 13.355 4.215 ;
      RECT  9.12 4.215 13.355 4.235 ;
      RECT  9.12 4.235 12.435 4.445 ;
      RECT  9.12 4.445 9.35 4.465 ;
      RECT  8.44 4.465 9.35 4.695 ;
      RECT  13.595 3.805 18.44 4.035 ;
      RECT  13.595 4.035 13.825 4.48 ;
      RECT  12.92 4.48 13.825 4.71 ;
      RECT  4.365 4.215 6.835 4.365 ;
      RECT  4.365 4.365 7.24 4.445 ;
      RECT  4.365 4.445 4.595 4.54 ;
      RECT  6.605 4.445 7.24 4.595 ;
      RECT  3.245 4.54 4.595 4.77 ;
      RECT  3.245 4.77 3.475 5.21 ;
      RECT  14.06 4.365 17.42 4.595 ;
      RECT  14.06 4.595 14.29 4.81 ;
      RECT  17.19 4.595 17.42 5.0 ;
      RECT  14.055 4.81 14.29 4.815 ;
      RECT  14.05 4.815 14.29 4.82 ;
      RECT  14.045 4.82 14.29 4.825 ;
      RECT  14.04 4.825 14.29 4.83 ;
      RECT  14.035 4.83 14.29 4.835 ;
      RECT  14.03 4.835 14.29 4.84 ;
      RECT  14.025 4.84 14.29 4.845 ;
      RECT  14.02 4.845 14.29 4.85 ;
      RECT  14.015 4.85 14.29 4.855 ;
      RECT  14.01 4.855 14.29 4.86 ;
      RECT  14.005 4.86 14.29 4.865 ;
      RECT  14.0 4.865 14.29 4.87 ;
      RECT  13.995 4.87 14.29 4.875 ;
      RECT  13.99 4.875 14.29 4.88 ;
      RECT  13.985 4.88 14.29 4.885 ;
      RECT  13.98 4.885 14.29 4.89 ;
      RECT  13.975 4.89 14.29 4.895 ;
      RECT  13.97 4.895 14.29 4.9 ;
      RECT  13.965 4.9 14.29 4.905 ;
      RECT  13.96 4.905 14.285 4.91 ;
      RECT  13.955 4.91 14.28 4.915 ;
      RECT  13.95 4.915 14.275 4.92 ;
      RECT  13.945 4.92 14.27 4.925 ;
      RECT  13.94 4.925 14.265 4.93 ;
      RECT  13.935 4.93 14.26 4.935 ;
      RECT  13.93 4.935 14.255 4.94 ;
      RECT  13.925 4.94 14.25 4.945 ;
      RECT  13.92 4.945 14.245 4.95 ;
      RECT  13.915 4.95 14.24 4.955 ;
      RECT  13.91 4.955 14.235 4.96 ;
      RECT  13.905 4.96 14.23 4.965 ;
      RECT  13.9 4.965 14.225 4.97 ;
      RECT  13.895 4.97 14.22 4.975 ;
      RECT  13.89 4.975 14.215 4.98 ;
      RECT  12.15 4.98 14.21 4.985 ;
      RECT  12.15 4.985 14.205 4.99 ;
      RECT  12.15 4.99 14.2 4.995 ;
      RECT  12.15 4.995 14.195 5.0 ;
      RECT  12.15 5.0 14.19 5.005 ;
      RECT  17.19 5.0 17.53 5.23 ;
      RECT  12.15 5.005 14.185 5.01 ;
      RECT  12.15 5.01 14.18 5.015 ;
      RECT  12.15 5.015 14.175 5.02 ;
      RECT  12.15 5.02 14.17 5.025 ;
      RECT  12.15 5.025 14.165 5.03 ;
      RECT  12.15 5.03 14.16 5.035 ;
      RECT  12.15 5.035 14.155 5.04 ;
      RECT  12.15 5.04 14.15 5.045 ;
      RECT  12.15 5.045 14.145 5.05 ;
      RECT  12.15 5.05 14.14 5.055 ;
      RECT  12.15 5.055 14.135 5.06 ;
      RECT  12.15 5.06 14.13 5.065 ;
      RECT  12.15 5.065 14.125 5.07 ;
      RECT  12.15 5.07 14.12 5.075 ;
      RECT  12.15 5.075 14.115 5.08 ;
      RECT  12.15 5.08 14.11 5.085 ;
      RECT  12.15 5.085 14.105 5.09 ;
      RECT  12.15 5.09 14.1 5.095 ;
      RECT  12.15 5.095 14.095 5.1 ;
      RECT  12.15 5.1 14.09 5.105 ;
      RECT  12.15 5.105 14.085 5.11 ;
      RECT  12.15 5.11 14.08 5.115 ;
      RECT  12.15 5.115 14.075 5.12 ;
      RECT  12.15 5.12 14.07 5.125 ;
      RECT  12.15 5.125 14.065 5.13 ;
      RECT  12.15 5.13 14.06 5.135 ;
      RECT  12.15 5.135 14.055 5.14 ;
      RECT  12.15 5.14 14.05 5.145 ;
      RECT  12.15 5.145 14.045 5.15 ;
      RECT  12.15 5.15 14.04 5.155 ;
      RECT  12.15 5.155 14.035 5.16 ;
      RECT  12.15 5.16 14.03 5.165 ;
      RECT  12.15 5.165 14.025 5.17 ;
      RECT  12.15 5.17 14.02 5.175 ;
      RECT  12.15 5.175 14.015 5.18 ;
      RECT  12.15 5.18 14.01 5.185 ;
      RECT  12.15 5.185 14.005 5.19 ;
      RECT  12.15 5.19 14.0 5.195 ;
      RECT  12.15 5.195 13.995 5.2 ;
      RECT  12.15 5.2 13.99 5.205 ;
      RECT  12.15 5.205 13.985 5.21 ;
      RECT  9.71 4.675 10.755 4.68 ;
      RECT  9.705 4.68 10.755 4.685 ;
      RECT  9.7 4.685 10.755 4.69 ;
      RECT  9.695 4.69 10.755 4.695 ;
      RECT  9.69 4.695 10.755 4.7 ;
      RECT  9.685 4.7 10.755 4.705 ;
      RECT  9.68 4.705 10.755 4.71 ;
      RECT  9.675 4.71 10.755 4.715 ;
      RECT  9.67 4.715 10.755 4.72 ;
      RECT  9.665 4.72 10.755 4.725 ;
      RECT  9.66 4.725 10.755 4.73 ;
      RECT  9.655 4.73 10.755 4.735 ;
      RECT  9.65 4.735 10.755 4.74 ;
      RECT  9.645 4.74 10.755 4.745 ;
      RECT  9.64 4.745 10.755 4.75 ;
      RECT  9.635 4.75 10.755 4.755 ;
      RECT  9.63 4.755 10.755 4.76 ;
      RECT  9.625 4.76 10.755 4.765 ;
      RECT  9.62 4.765 10.755 4.77 ;
      RECT  9.615 4.77 10.755 4.775 ;
      RECT  9.61 4.775 10.755 4.78 ;
      RECT  9.605 4.78 10.755 4.785 ;
      RECT  9.6 4.785 10.755 4.79 ;
      RECT  9.595 4.79 10.755 4.795 ;
      RECT  9.59 4.795 10.755 4.8 ;
      RECT  9.585 4.8 10.755 4.805 ;
      RECT  9.58 4.805 10.755 4.81 ;
      RECT  9.575 4.81 10.755 4.815 ;
      RECT  9.57 4.815 10.755 4.82 ;
      RECT  9.565 4.82 10.755 4.825 ;
      RECT  9.56 4.825 10.755 4.83 ;
      RECT  9.555 4.83 10.755 4.835 ;
      RECT  9.55 4.835 10.755 4.84 ;
      RECT  9.545 4.84 10.755 4.845 ;
      RECT  9.54 4.845 10.755 4.85 ;
      RECT  9.535 4.85 10.755 4.855 ;
      RECT  9.53 4.855 10.755 4.86 ;
      RECT  9.525 4.86 10.755 4.865 ;
      RECT  9.52 4.865 10.755 4.87 ;
      RECT  9.515 4.87 10.755 4.875 ;
      RECT  9.51 4.875 10.755 4.88 ;
      RECT  9.505 4.88 10.755 4.885 ;
      RECT  9.5 4.885 10.755 4.89 ;
      RECT  9.495 4.89 10.755 4.895 ;
      RECT  9.49 4.895 10.755 4.9 ;
      RECT  9.485 4.9 10.755 4.905 ;
      RECT  9.48 4.905 9.805 4.91 ;
      RECT  10.525 4.905 10.755 5.0 ;
      RECT  9.475 4.91 9.8 4.915 ;
      RECT  9.47 4.915 9.795 4.92 ;
      RECT  9.465 4.92 9.79 4.925 ;
      RECT  9.46 4.925 9.785 4.93 ;
      RECT  9.455 4.93 9.78 4.935 ;
      RECT  9.45 4.935 9.775 4.94 ;
      RECT  9.445 4.94 9.77 4.945 ;
      RECT  9.44 4.945 9.765 4.95 ;
      RECT  9.435 4.95 9.76 4.955 ;
      RECT  9.43 4.955 9.755 4.96 ;
      RECT  9.425 4.96 9.75 4.965 ;
      RECT  9.42 4.965 9.745 4.97 ;
      RECT  9.415 4.97 9.74 4.975 ;
      RECT  9.41 4.975 9.735 4.98 ;
      RECT  9.405 4.98 9.73 4.985 ;
      RECT  9.4 4.985 9.725 4.99 ;
      RECT  9.395 4.99 9.72 4.995 ;
      RECT  9.39 4.995 9.715 5.0 ;
      RECT  8.23 5.0 9.71 5.005 ;
      RECT  10.525 5.0 11.91 5.23 ;
      RECT  8.23 5.005 9.705 5.01 ;
      RECT  8.23 5.01 9.7 5.015 ;
      RECT  8.23 5.015 9.695 5.02 ;
      RECT  8.23 5.02 9.69 5.025 ;
      RECT  8.23 5.025 9.685 5.03 ;
      RECT  8.23 5.03 9.68 5.035 ;
      RECT  8.23 5.035 9.675 5.04 ;
      RECT  8.23 5.04 9.67 5.045 ;
      RECT  8.23 5.045 9.665 5.05 ;
      RECT  8.23 5.05 9.66 5.055 ;
      RECT  8.23 5.055 9.655 5.06 ;
      RECT  8.23 5.06 9.65 5.065 ;
      RECT  8.23 5.065 9.645 5.07 ;
      RECT  8.23 5.07 9.64 5.075 ;
      RECT  8.23 5.075 9.635 5.08 ;
      RECT  8.23 5.08 9.63 5.085 ;
      RECT  8.23 5.085 9.625 5.09 ;
      RECT  8.23 5.09 9.62 5.095 ;
      RECT  8.23 5.095 9.615 5.1 ;
      RECT  8.23 5.1 9.61 5.105 ;
      RECT  8.23 5.105 9.605 5.11 ;
      RECT  8.23 5.11 9.6 5.115 ;
      RECT  8.23 5.115 9.595 5.12 ;
      RECT  8.23 5.12 9.59 5.125 ;
      RECT  8.23 5.125 9.585 5.13 ;
      RECT  8.23 5.13 9.58 5.135 ;
      RECT  8.23 5.135 9.575 5.14 ;
      RECT  8.23 5.14 9.57 5.145 ;
      RECT  8.23 5.145 9.565 5.15 ;
      RECT  8.23 5.15 9.56 5.155 ;
      RECT  8.23 5.155 9.555 5.16 ;
      RECT  8.23 5.16 9.55 5.165 ;
      RECT  8.23 5.165 9.545 5.17 ;
      RECT  8.23 5.17 9.54 5.175 ;
      RECT  8.23 5.175 9.535 5.18 ;
      RECT  8.23 5.18 9.53 5.185 ;
      RECT  8.23 5.185 9.525 5.19 ;
      RECT  8.23 5.19 9.52 5.195 ;
      RECT  8.23 5.195 9.515 5.2 ;
      RECT  8.23 5.2 9.51 5.205 ;
      RECT  8.23 5.205 9.505 5.21 ;
      RECT  8.23 5.21 9.5 5.215 ;
      RECT  8.23 5.215 9.495 5.22 ;
      RECT  8.23 5.22 9.49 5.225 ;
      RECT  8.23 5.225 9.485 5.23 ;
      LAYER METAL2 ;
      RECT  8.77 2.66 10.83 2.94 ;
      LAYER VIA12 ;
      RECT  8.83 2.67 9.09 2.93 ;
      RECT  10.51 2.67 10.77 2.93 ;
  END
END MDN_FSDNRBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNRBQ_4
#      Description : D-Flip Flop w/scan, neg-edge triggered, lo-async-clear, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNRBQ_4
  CLASS CORE ;
  FOREIGN MDN_FSDNRBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 24.64 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 1.565 2.94 2.69 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.64 1.565 22.92 1.795 ;
      RECT  22.285 1.795 22.515 3.245 ;
      RECT  19.64 3.245 22.92 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.98 2.125 16.38 2.355 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.81 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  20.72 5.46 21.395 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  16.63 5.135 16.97 5.46 ;
      RECT  16.24 5.46 17.36 5.74 ;
      RECT  14.39 5.135 14.73 5.46 ;
      RECT  14.0 5.46 15.12 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 11.37 5.74 ;
      RECT  5.43 5.135 5.77 5.46 ;
      RECT  5.04 5.46 6.16 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 24.64 5.74 ;
      LAYER VIA12 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  24.23 5.47 24.49 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 24.81 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  15.12 -0.14 16.24 0.14 ;
      RECT  15.565 0.14 15.795 1.005 ;
      RECT  15.16 1.005 16.2 1.235 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.6 ;
      RECT  3.805 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.6 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 24.64 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  22.55 -0.13 22.81 0.13 ;
      RECT  23.11 -0.13 23.37 0.13 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  10.425 0.37 13.05 0.6 ;
      RECT  10.425 0.6 10.655 0.83 ;
      RECT  5.98 0.37 9.635 0.6 ;
      RECT  5.98 0.6 6.21 0.83 ;
      RECT  9.405 0.6 9.635 0.83 ;
      RECT  4.715 0.83 6.21 1.06 ;
      RECT  9.405 0.83 10.655 1.06 ;
      RECT  4.715 1.06 4.945 1.29 ;
      RECT  21.67 0.37 23.13 0.6 ;
      RECT  6.44 0.83 8.78 1.06 ;
      RECT  8.44 1.06 8.78 1.12 ;
      RECT  6.44 1.06 6.67 1.29 ;
      RECT  5.485 1.29 6.67 1.52 ;
      RECT  5.485 1.52 5.715 1.565 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  3.245 1.565 5.715 1.795 ;
      RECT  10.885 0.83 13.96 1.06 ;
      RECT  13.62 1.06 13.96 1.12 ;
      RECT  10.885 1.06 11.115 1.29 ;
      RECT  8.945 1.29 11.115 1.295 ;
      RECT  8.94 1.295 11.115 1.3 ;
      RECT  8.935 1.3 11.115 1.305 ;
      RECT  8.93 1.305 11.115 1.31 ;
      RECT  8.925 1.31 11.115 1.315 ;
      RECT  8.92 1.315 11.115 1.32 ;
      RECT  8.915 1.32 11.115 1.325 ;
      RECT  8.91 1.325 11.115 1.33 ;
      RECT  8.905 1.33 11.115 1.335 ;
      RECT  8.9 1.335 11.115 1.34 ;
      RECT  8.895 1.34 11.115 1.345 ;
      RECT  8.89 1.345 11.115 1.35 ;
      RECT  6.9 1.29 8.27 1.35 ;
      RECT  6.9 1.35 11.115 1.52 ;
      RECT  8.115 1.52 9.04 1.525 ;
      RECT  8.115 1.525 9.035 1.53 ;
      RECT  8.115 1.53 9.03 1.535 ;
      RECT  8.115 1.535 9.025 1.54 ;
      RECT  8.115 1.54 9.02 1.545 ;
      RECT  8.115 1.545 9.015 1.55 ;
      RECT  8.115 1.55 9.01 1.555 ;
      RECT  8.115 1.555 9.005 1.56 ;
      RECT  8.115 1.56 9.0 1.565 ;
      RECT  8.115 1.565 8.995 1.57 ;
      RECT  8.115 1.57 8.99 1.575 ;
      RECT  8.115 1.575 8.985 1.58 ;
      RECT  16.685 1.005 18.44 1.235 ;
      RECT  16.685 1.235 16.915 1.565 ;
      RECT  11.38 1.29 13.465 1.295 ;
      RECT  11.38 1.295 13.47 1.3 ;
      RECT  11.38 1.3 13.475 1.305 ;
      RECT  11.38 1.305 13.48 1.31 ;
      RECT  11.38 1.31 13.485 1.315 ;
      RECT  11.38 1.315 13.49 1.32 ;
      RECT  11.38 1.32 13.495 1.325 ;
      RECT  11.38 1.325 13.5 1.33 ;
      RECT  11.38 1.33 13.505 1.335 ;
      RECT  11.38 1.335 13.51 1.34 ;
      RECT  11.38 1.34 13.515 1.345 ;
      RECT  11.38 1.345 13.52 1.35 ;
      RECT  11.38 1.35 13.525 1.355 ;
      RECT  11.38 1.355 13.53 1.36 ;
      RECT  11.38 1.36 13.535 1.365 ;
      RECT  11.38 1.365 13.54 1.37 ;
      RECT  11.38 1.37 13.545 1.375 ;
      RECT  11.38 1.375 13.55 1.38 ;
      RECT  11.38 1.38 13.555 1.385 ;
      RECT  11.38 1.385 13.56 1.39 ;
      RECT  11.38 1.39 13.565 1.395 ;
      RECT  11.38 1.395 13.57 1.4 ;
      RECT  11.38 1.4 13.575 1.405 ;
      RECT  11.38 1.405 13.58 1.41 ;
      RECT  11.38 1.41 13.585 1.415 ;
      RECT  11.38 1.415 13.59 1.42 ;
      RECT  11.38 1.42 13.595 1.425 ;
      RECT  11.38 1.425 13.6 1.43 ;
      RECT  11.38 1.43 13.605 1.435 ;
      RECT  11.38 1.435 13.61 1.44 ;
      RECT  11.38 1.44 13.615 1.445 ;
      RECT  11.38 1.445 13.62 1.45 ;
      RECT  11.38 1.45 13.625 1.455 ;
      RECT  11.38 1.455 13.63 1.46 ;
      RECT  11.38 1.46 13.635 1.465 ;
      RECT  11.38 1.465 13.64 1.47 ;
      RECT  11.38 1.47 13.645 1.475 ;
      RECT  11.38 1.475 13.65 1.48 ;
      RECT  11.38 1.48 13.655 1.485 ;
      RECT  11.38 1.485 13.66 1.49 ;
      RECT  11.38 1.49 13.665 1.495 ;
      RECT  11.38 1.495 13.67 1.5 ;
      RECT  11.38 1.5 13.675 1.505 ;
      RECT  11.38 1.505 13.68 1.51 ;
      RECT  11.38 1.51 13.685 1.515 ;
      RECT  11.38 1.515 13.69 1.52 ;
      RECT  13.36 1.52 13.695 1.525 ;
      RECT  13.365 1.525 13.7 1.53 ;
      RECT  13.37 1.53 13.705 1.535 ;
      RECT  13.375 1.535 13.71 1.54 ;
      RECT  13.38 1.54 13.715 1.545 ;
      RECT  13.385 1.545 13.72 1.55 ;
      RECT  13.39 1.55 13.725 1.555 ;
      RECT  13.395 1.555 13.73 1.56 ;
      RECT  13.4 1.56 13.735 1.565 ;
      RECT  13.405 1.565 16.915 1.57 ;
      RECT  13.41 1.57 16.915 1.575 ;
      RECT  13.415 1.575 16.915 1.58 ;
      RECT  13.42 1.58 16.915 1.585 ;
      RECT  13.425 1.585 16.915 1.59 ;
      RECT  13.43 1.59 16.915 1.595 ;
      RECT  13.435 1.595 16.915 1.6 ;
      RECT  13.44 1.6 16.915 1.605 ;
      RECT  13.445 1.605 16.915 1.61 ;
      RECT  13.45 1.61 16.915 1.615 ;
      RECT  13.455 1.615 16.915 1.62 ;
      RECT  13.46 1.62 16.915 1.625 ;
      RECT  13.465 1.625 16.915 1.63 ;
      RECT  13.47 1.63 16.915 1.635 ;
      RECT  13.475 1.635 16.915 1.64 ;
      RECT  13.48 1.64 16.915 1.645 ;
      RECT  13.485 1.645 16.915 1.65 ;
      RECT  13.49 1.65 16.915 1.655 ;
      RECT  13.495 1.655 16.915 1.66 ;
      RECT  13.5 1.66 16.915 1.665 ;
      RECT  13.505 1.665 16.915 1.67 ;
      RECT  13.51 1.67 16.915 1.675 ;
      RECT  13.515 1.675 16.915 1.68 ;
      RECT  13.52 1.68 16.915 1.685 ;
      RECT  13.525 1.685 16.915 1.69 ;
      RECT  13.53 1.69 16.915 1.695 ;
      RECT  13.535 1.695 16.915 1.7 ;
      RECT  13.54 1.7 16.915 1.705 ;
      RECT  13.545 1.705 16.915 1.71 ;
      RECT  13.55 1.71 16.915 1.715 ;
      RECT  13.555 1.715 16.915 1.72 ;
      RECT  13.56 1.72 16.915 1.725 ;
      RECT  13.565 1.725 16.915 1.73 ;
      RECT  13.57 1.73 16.915 1.735 ;
      RECT  13.575 1.735 16.915 1.74 ;
      RECT  13.58 1.74 16.915 1.745 ;
      RECT  13.585 1.745 16.915 1.75 ;
      RECT  13.59 1.75 16.915 1.755 ;
      RECT  13.595 1.755 16.915 1.76 ;
      RECT  13.6 1.76 16.915 1.765 ;
      RECT  13.605 1.765 16.915 1.77 ;
      RECT  13.61 1.77 16.915 1.775 ;
      RECT  13.615 1.775 16.915 1.78 ;
      RECT  13.62 1.78 16.915 1.785 ;
      RECT  13.625 1.785 16.915 1.79 ;
      RECT  13.63 1.79 16.915 1.795 ;
      RECT  17.4 1.565 18.595 1.795 ;
      RECT  18.365 1.795 18.595 2.405 ;
      RECT  18.365 2.405 21.825 2.635 ;
      RECT  18.365 2.635 18.595 3.245 ;
      RECT  15.86 3.245 18.595 3.475 ;
      RECT  7.62 1.75 7.96 1.82 ;
      RECT  7.62 1.82 8.865 2.05 ;
      RECT  8.635 2.05 8.865 2.66 ;
      RECT  8.635 2.66 9.15 2.8 ;
      RECT  7.725 2.8 9.15 2.94 ;
      RECT  7.725 2.94 8.87 3.03 ;
      RECT  7.725 3.03 7.955 3.315 ;
      RECT  6.2 1.75 6.835 1.98 ;
      RECT  6.605 1.98 6.835 2.34 ;
      RECT  6.605 2.34 8.405 2.57 ;
      RECT  6.605 2.57 6.835 3.245 ;
      RECT  6.2 3.245 6.835 3.475 ;
      RECT  9.14 1.75 10.195 1.98 ;
      RECT  9.965 1.98 10.195 3.72 ;
      RECT  8.655 3.72 10.195 3.95 ;
      RECT  8.655 3.95 8.885 4.02 ;
      RECT  7.725 4.02 8.885 4.25 ;
      RECT  7.725 4.25 7.955 4.925 ;
      RECT  4.925 4.675 6.275 4.905 ;
      RECT  6.045 4.905 6.275 4.925 ;
      RECT  4.925 4.905 5.155 5.0 ;
      RECT  6.045 4.925 7.955 5.155 ;
      RECT  3.75 5.0 5.155 5.23 ;
      RECT  12.15 1.75 12.49 1.98 ;
      RECT  12.205 1.98 12.435 3.315 ;
      RECT  12.765 1.75 13.26 1.98 ;
      RECT  12.765 1.98 12.995 2.685 ;
      RECT  12.665 2.685 14.115 2.915 ;
      RECT  13.885 2.35 14.115 2.685 ;
      RECT  12.665 2.915 12.895 3.545 ;
      RECT  10.68 1.75 11.315 1.98 ;
      RECT  11.085 1.98 11.315 3.545 ;
      RECT  10.68 3.545 12.895 3.775 ;
      RECT  5.485 2.41 6.33 2.64 ;
      RECT  5.485 2.64 5.715 3.245 ;
      RECT  4.66 3.245 5.715 3.475 ;
      RECT  10.47 2.28 10.81 2.66 ;
      RECT  10.43 2.66 10.81 2.94 ;
      RECT  9.405 2.35 9.635 3.26 ;
      RECT  8.195 3.26 9.635 3.49 ;
      RECT  8.195 3.49 8.425 3.56 ;
      RECT  7.165 3.56 8.425 3.755 ;
      RECT  3.805 3.755 8.425 3.79 ;
      RECT  3.805 3.79 7.395 3.985 ;
      RECT  3.805 3.985 4.035 4.08 ;
      RECT  2.685 4.08 4.035 4.31 ;
      RECT  2.685 4.31 2.915 4.37 ;
      RECT  1.51 4.37 2.915 4.6 ;
      RECT  1.51 4.6 1.74 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  1.72 3.16 2.76 3.39 ;
      RECT  3.245 3.245 4.3 3.475 ;
      RECT  3.245 3.475 3.475 3.62 ;
      RECT  2.115 3.62 3.475 3.805 ;
      RECT  0.18 3.805 3.475 3.85 ;
      RECT  0.18 3.85 2.35 4.035 ;
      RECT  13.125 3.245 15.5 3.475 ;
      RECT  13.125 3.475 13.355 4.02 ;
      RECT  12.205 4.02 13.355 4.215 ;
      RECT  9.115 4.215 13.355 4.25 ;
      RECT  9.115 4.25 12.435 4.445 ;
      RECT  9.115 4.445 9.345 4.48 ;
      RECT  8.44 4.48 9.345 4.71 ;
      RECT  13.585 3.805 18.44 4.035 ;
      RECT  13.585 4.035 13.815 4.48 ;
      RECT  12.92 4.48 13.815 4.71 ;
      RECT  4.365 4.215 7.245 4.445 ;
      RECT  4.365 4.445 4.595 4.54 ;
      RECT  3.245 4.54 4.595 4.77 ;
      RECT  3.245 4.77 3.475 5.21 ;
      RECT  14.075 4.37 17.43 4.6 ;
      RECT  14.075 4.6 14.305 4.795 ;
      RECT  17.2 4.6 17.43 5.0 ;
      RECT  14.07 4.795 14.305 4.8 ;
      RECT  14.065 4.8 14.305 4.805 ;
      RECT  14.06 4.805 14.305 4.81 ;
      RECT  14.055 4.81 14.305 4.815 ;
      RECT  14.05 4.815 14.305 4.82 ;
      RECT  14.045 4.82 14.305 4.825 ;
      RECT  14.04 4.825 14.305 4.83 ;
      RECT  14.035 4.83 14.305 4.835 ;
      RECT  14.03 4.835 14.305 4.84 ;
      RECT  14.025 4.84 14.305 4.845 ;
      RECT  14.02 4.845 14.305 4.85 ;
      RECT  14.015 4.85 14.305 4.855 ;
      RECT  14.01 4.855 14.305 4.86 ;
      RECT  14.005 4.86 14.305 4.865 ;
      RECT  14.0 4.865 14.305 4.87 ;
      RECT  13.995 4.87 14.305 4.875 ;
      RECT  13.99 4.875 14.305 4.88 ;
      RECT  13.985 4.88 14.305 4.885 ;
      RECT  13.98 4.885 14.305 4.89 ;
      RECT  13.975 4.89 14.3 4.895 ;
      RECT  13.97 4.895 14.295 4.9 ;
      RECT  13.965 4.9 14.29 4.905 ;
      RECT  13.96 4.905 14.285 4.91 ;
      RECT  13.955 4.91 14.28 4.915 ;
      RECT  13.95 4.915 14.275 4.92 ;
      RECT  13.945 4.92 14.27 4.925 ;
      RECT  13.94 4.925 14.265 4.93 ;
      RECT  13.935 4.93 14.26 4.935 ;
      RECT  13.93 4.935 14.255 4.94 ;
      RECT  13.925 4.94 14.25 4.945 ;
      RECT  13.92 4.945 14.245 4.95 ;
      RECT  13.915 4.95 14.24 4.955 ;
      RECT  13.91 4.955 14.235 4.96 ;
      RECT  13.905 4.96 14.23 4.965 ;
      RECT  13.9 4.965 14.225 4.97 ;
      RECT  13.895 4.97 14.22 4.975 ;
      RECT  13.89 4.975 14.215 4.98 ;
      RECT  12.15 4.98 14.21 4.985 ;
      RECT  12.15 4.985 14.205 4.99 ;
      RECT  12.15 4.99 14.2 4.995 ;
      RECT  12.15 4.995 14.195 5.0 ;
      RECT  12.15 5.0 14.19 5.005 ;
      RECT  17.2 5.0 17.54 5.23 ;
      RECT  12.15 5.005 14.185 5.01 ;
      RECT  12.15 5.01 14.18 5.015 ;
      RECT  12.15 5.015 14.175 5.02 ;
      RECT  12.15 5.02 14.17 5.025 ;
      RECT  12.15 5.025 14.165 5.03 ;
      RECT  12.15 5.03 14.16 5.035 ;
      RECT  12.15 5.035 14.155 5.04 ;
      RECT  12.15 5.04 14.15 5.045 ;
      RECT  12.15 5.045 14.145 5.05 ;
      RECT  12.15 5.05 14.14 5.055 ;
      RECT  12.15 5.055 14.135 5.06 ;
      RECT  12.15 5.06 14.13 5.065 ;
      RECT  12.15 5.065 14.125 5.07 ;
      RECT  12.15 5.07 14.12 5.075 ;
      RECT  12.15 5.075 14.115 5.08 ;
      RECT  12.15 5.08 14.11 5.085 ;
      RECT  12.15 5.085 14.105 5.09 ;
      RECT  12.15 5.09 14.1 5.095 ;
      RECT  12.15 5.095 14.095 5.1 ;
      RECT  12.15 5.1 14.09 5.105 ;
      RECT  12.15 5.105 14.085 5.11 ;
      RECT  12.15 5.11 14.08 5.115 ;
      RECT  12.15 5.115 14.075 5.12 ;
      RECT  12.15 5.12 14.07 5.125 ;
      RECT  12.15 5.125 14.065 5.13 ;
      RECT  12.15 5.13 14.06 5.135 ;
      RECT  12.15 5.135 14.055 5.14 ;
      RECT  12.15 5.14 14.05 5.145 ;
      RECT  12.15 5.145 14.045 5.15 ;
      RECT  12.15 5.15 14.04 5.155 ;
      RECT  12.15 5.155 14.035 5.16 ;
      RECT  12.15 5.16 14.03 5.165 ;
      RECT  12.15 5.165 14.025 5.17 ;
      RECT  12.15 5.17 14.02 5.175 ;
      RECT  12.15 5.175 14.015 5.18 ;
      RECT  12.15 5.18 14.01 5.185 ;
      RECT  12.15 5.185 14.005 5.19 ;
      RECT  12.15 5.19 14.0 5.195 ;
      RECT  12.15 5.195 13.995 5.2 ;
      RECT  12.15 5.2 13.99 5.205 ;
      RECT  12.15 5.205 13.985 5.21 ;
      RECT  9.71 4.675 10.755 4.68 ;
      RECT  9.705 4.68 10.755 4.685 ;
      RECT  9.7 4.685 10.755 4.69 ;
      RECT  9.695 4.69 10.755 4.695 ;
      RECT  9.69 4.695 10.755 4.7 ;
      RECT  9.685 4.7 10.755 4.705 ;
      RECT  9.68 4.705 10.755 4.71 ;
      RECT  9.675 4.71 10.755 4.715 ;
      RECT  9.67 4.715 10.755 4.72 ;
      RECT  9.665 4.72 10.755 4.725 ;
      RECT  9.66 4.725 10.755 4.73 ;
      RECT  9.655 4.73 10.755 4.735 ;
      RECT  9.65 4.735 10.755 4.74 ;
      RECT  9.645 4.74 10.755 4.745 ;
      RECT  9.64 4.745 10.755 4.75 ;
      RECT  9.635 4.75 10.755 4.755 ;
      RECT  9.63 4.755 10.755 4.76 ;
      RECT  9.625 4.76 10.755 4.765 ;
      RECT  9.62 4.765 10.755 4.77 ;
      RECT  9.615 4.77 10.755 4.775 ;
      RECT  9.61 4.775 10.755 4.78 ;
      RECT  9.605 4.78 10.755 4.785 ;
      RECT  9.6 4.785 10.755 4.79 ;
      RECT  9.595 4.79 10.755 4.795 ;
      RECT  9.59 4.795 10.755 4.8 ;
      RECT  9.585 4.8 10.755 4.805 ;
      RECT  9.58 4.805 10.755 4.81 ;
      RECT  9.575 4.81 10.755 4.815 ;
      RECT  9.57 4.815 10.755 4.82 ;
      RECT  9.565 4.82 10.755 4.825 ;
      RECT  9.56 4.825 10.755 4.83 ;
      RECT  9.555 4.83 10.755 4.835 ;
      RECT  9.55 4.835 10.755 4.84 ;
      RECT  9.545 4.84 10.755 4.845 ;
      RECT  9.54 4.845 10.755 4.85 ;
      RECT  9.535 4.85 10.755 4.855 ;
      RECT  9.53 4.855 10.755 4.86 ;
      RECT  9.525 4.86 10.755 4.865 ;
      RECT  9.52 4.865 10.755 4.87 ;
      RECT  9.515 4.87 10.755 4.875 ;
      RECT  9.51 4.875 10.755 4.88 ;
      RECT  9.505 4.88 10.755 4.885 ;
      RECT  9.5 4.885 10.755 4.89 ;
      RECT  9.495 4.89 10.755 4.895 ;
      RECT  9.49 4.895 10.755 4.9 ;
      RECT  9.485 4.9 10.755 4.905 ;
      RECT  9.48 4.905 9.805 4.91 ;
      RECT  10.525 4.905 10.755 5.0 ;
      RECT  9.475 4.91 9.8 4.915 ;
      RECT  9.47 4.915 9.795 4.92 ;
      RECT  9.465 4.92 9.79 4.925 ;
      RECT  9.46 4.925 9.785 4.93 ;
      RECT  9.455 4.93 9.78 4.935 ;
      RECT  9.45 4.935 9.775 4.94 ;
      RECT  9.445 4.94 9.77 4.945 ;
      RECT  9.44 4.945 9.765 4.95 ;
      RECT  9.435 4.95 9.76 4.955 ;
      RECT  9.43 4.955 9.755 4.96 ;
      RECT  9.425 4.96 9.75 4.965 ;
      RECT  9.42 4.965 9.745 4.97 ;
      RECT  9.415 4.97 9.74 4.975 ;
      RECT  9.41 4.975 9.735 4.98 ;
      RECT  9.405 4.98 9.73 4.985 ;
      RECT  9.4 4.985 9.725 4.99 ;
      RECT  9.395 4.99 9.72 4.995 ;
      RECT  9.39 4.995 9.715 5.0 ;
      RECT  8.23 5.0 9.71 5.005 ;
      RECT  10.525 5.0 11.91 5.23 ;
      RECT  8.23 5.005 9.705 5.01 ;
      RECT  8.23 5.01 9.7 5.015 ;
      RECT  8.23 5.015 9.695 5.02 ;
      RECT  8.23 5.02 9.69 5.025 ;
      RECT  8.23 5.025 9.685 5.03 ;
      RECT  8.23 5.03 9.68 5.035 ;
      RECT  8.23 5.035 9.675 5.04 ;
      RECT  8.23 5.04 9.67 5.045 ;
      RECT  8.23 5.045 9.665 5.05 ;
      RECT  8.23 5.05 9.66 5.055 ;
      RECT  8.23 5.055 9.655 5.06 ;
      RECT  8.23 5.06 9.65 5.065 ;
      RECT  8.23 5.065 9.645 5.07 ;
      RECT  8.23 5.07 9.64 5.075 ;
      RECT  8.23 5.075 9.635 5.08 ;
      RECT  8.23 5.08 9.63 5.085 ;
      RECT  8.23 5.085 9.625 5.09 ;
      RECT  8.23 5.09 9.62 5.095 ;
      RECT  8.23 5.095 9.615 5.1 ;
      RECT  8.23 5.1 9.61 5.105 ;
      RECT  8.23 5.105 9.605 5.11 ;
      RECT  8.23 5.11 9.6 5.115 ;
      RECT  8.23 5.115 9.595 5.12 ;
      RECT  8.23 5.12 9.59 5.125 ;
      RECT  8.23 5.125 9.585 5.13 ;
      RECT  8.23 5.13 9.58 5.135 ;
      RECT  8.23 5.135 9.575 5.14 ;
      RECT  8.23 5.14 9.57 5.145 ;
      RECT  8.23 5.145 9.565 5.15 ;
      RECT  8.23 5.15 9.56 5.155 ;
      RECT  8.23 5.155 9.555 5.16 ;
      RECT  8.23 5.16 9.55 5.165 ;
      RECT  8.23 5.165 9.545 5.17 ;
      RECT  8.23 5.17 9.54 5.175 ;
      RECT  8.23 5.175 9.535 5.18 ;
      RECT  8.23 5.18 9.53 5.185 ;
      RECT  8.23 5.185 9.525 5.19 ;
      RECT  8.23 5.19 9.52 5.195 ;
      RECT  8.23 5.195 9.515 5.2 ;
      RECT  8.23 5.2 9.51 5.205 ;
      RECT  8.23 5.205 9.505 5.21 ;
      RECT  8.23 5.21 9.5 5.215 ;
      RECT  8.23 5.215 9.495 5.22 ;
      RECT  8.23 5.22 9.49 5.225 ;
      RECT  8.23 5.225 9.485 5.23 ;
      LAYER METAL2 ;
      RECT  8.77 2.66 10.81 2.94 ;
      LAYER VIA12 ;
      RECT  8.83 2.67 9.09 2.93 ;
      RECT  10.49 2.67 10.75 2.93 ;
  END
END MDN_FSDNRBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNRBSBQ_1
#      Description : D-Flip Flop w/scan, neg-edge triggered, lo-async-clear/set, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNRBSBQ_1
  CLASS CORE ;
  FOREIGN MDN_FSDNRBSBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 8.54 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  2.42 3.245 2.915 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.325 2.125 16.38 2.355 ;
      RECT  13.325 2.355 13.555 2.375 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  13.25 2.375 13.555 2.405 ;
      RECT  12.71 2.405 13.555 2.635 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.95 0.37 15.49 0.445 ;
      RECT  14.95 0.445 21.7 0.675 ;
      RECT  21.47 0.675 21.7 1.565 ;
      RECT  21.47 1.565 21.98 1.795 ;
      RECT  21.7 1.795 21.98 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 2.35 4.035 2.66 ;
      RECT  3.245 2.66 4.035 2.94 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.94 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  16.685 5.08 16.915 5.46 ;
      RECT  16.24 5.46 17.36 5.74 ;
      RECT  14.445 5.08 14.675 5.46 ;
      RECT  14.0 5.46 15.12 5.74 ;
      RECT  12.205 5.08 12.435 5.46 ;
      RECT  11.03 5.46 12.88 5.74 ;
      RECT  6.2 4.365 7.955 4.595 ;
      RECT  7.725 4.595 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.84 -0.14 22.57 0.14 ;
      RECT  21.935 0.14 22.165 1.175 ;
      RECT  14.0 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 1.005 ;
      RECT  12.92 1.005 16.2 1.235 ;
      RECT  11.03 -0.14 11.76 0.14 ;
      RECT  5.04 -0.14 6.16 0.14 ;
      RECT  5.43 0.14 5.77 0.465 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.52 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  13.83 0.37 14.17 0.445 ;
      RECT  12.205 0.445 14.17 0.675 ;
      RECT  12.205 0.675 12.435 1.48 ;
      RECT  11.085 1.48 12.435 1.565 ;
      RECT  9.91 1.565 12.435 1.71 ;
      RECT  9.91 1.71 11.315 1.795 ;
      RECT  11.085 1.795 11.315 3.03 ;
      RECT  9.91 3.03 11.315 3.26 ;
      RECT  1.465 0.37 1.85 0.6 ;
      RECT  1.465 0.6 1.695 0.98 ;
      RECT  1.315 0.98 1.695 1.005 ;
      RECT  0.18 1.005 1.695 1.235 ;
      RECT  1.315 1.235 1.695 1.26 ;
      RECT  6.045 0.37 9.69 0.6 ;
      RECT  6.045 0.6 6.275 0.695 ;
      RECT  3.805 0.695 6.275 0.925 ;
      RECT  3.805 0.925 4.035 1.005 ;
      RECT  1.925 1.005 4.035 1.235 ;
      RECT  1.925 1.235 2.155 1.565 ;
      RECT  1.565 1.565 2.155 1.795 ;
      RECT  1.565 1.795 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  10.185 0.37 10.81 0.6 ;
      RECT  10.185 0.6 10.415 0.98 ;
      RECT  9.89 0.98 10.415 1.26 ;
      RECT  6.605 1.005 8.78 1.155 ;
      RECT  4.66 1.155 8.78 1.235 ;
      RECT  4.66 1.235 6.835 1.385 ;
      RECT  18.1 0.945 20.625 1.175 ;
      RECT  20.395 1.175 20.625 1.285 ;
      RECT  10.68 1.005 11.72 1.235 ;
      RECT  20.855 0.98 21.235 1.26 ;
      RECT  20.855 1.26 21.085 1.565 ;
      RECT  20.605 1.565 21.085 1.795 ;
      RECT  20.605 1.795 20.835 2.39 ;
      RECT  19.655 2.39 20.835 2.62 ;
      RECT  18.365 1.405 19.21 1.635 ;
      RECT  18.365 1.635 18.595 2.335 ;
      RECT  17.19 2.335 18.595 2.565 ;
      RECT  18.365 2.565 18.595 3.24 ;
      RECT  18.365 3.24 19.16 3.47 ;
      RECT  7.67 1.565 9.51 1.795 ;
      RECT  12.765 1.565 13.96 1.795 ;
      RECT  12.765 1.795 12.995 1.94 ;
      RECT  11.645 1.94 12.995 2.17 ;
      RECT  11.645 2.17 11.875 3.03 ;
      RECT  11.645 3.03 13.96 3.26 ;
      RECT  16.685 1.565 17.74 1.795 ;
      RECT  16.685 1.795 16.915 3.24 ;
      RECT  15.565 3.24 17.74 3.47 ;
      RECT  15.565 3.47 15.795 3.49 ;
      RECT  4.925 3.245 9.075 3.475 ;
      RECT  8.845 3.475 9.075 3.49 ;
      RECT  4.925 3.475 5.155 3.805 ;
      RECT  8.845 3.49 15.795 3.72 ;
      RECT  3.805 3.805 5.155 4.035 ;
      RECT  3.805 4.035 4.035 4.365 ;
      RECT  2.74 4.365 4.035 4.595 ;
      RECT  2.74 4.595 2.97 5.0 ;
      RECT  2.63 5.0 2.97 5.23 ;
      RECT  6.2 1.62 7.24 1.85 ;
      RECT  19.64 1.75 19.98 1.865 ;
      RECT  18.925 1.865 19.98 2.095 ;
      RECT  18.925 2.095 19.155 2.555 ;
      RECT  18.925 2.555 19.16 2.56 ;
      RECT  18.925 2.56 19.165 2.565 ;
      RECT  18.925 2.565 19.17 2.57 ;
      RECT  18.925 2.57 19.175 2.575 ;
      RECT  18.925 2.575 19.18 2.58 ;
      RECT  18.925 2.58 19.185 2.585 ;
      RECT  18.925 2.585 19.19 2.59 ;
      RECT  18.925 2.59 19.195 2.595 ;
      RECT  18.925 2.595 19.2 2.6 ;
      RECT  18.925 2.6 19.205 2.605 ;
      RECT  18.925 2.605 19.21 2.61 ;
      RECT  18.925 2.61 19.215 2.615 ;
      RECT  18.925 2.615 19.22 2.62 ;
      RECT  18.925 2.62 19.225 2.625 ;
      RECT  18.925 2.625 19.23 2.63 ;
      RECT  18.925 2.63 19.235 2.635 ;
      RECT  18.925 2.635 19.24 2.64 ;
      RECT  18.925 2.64 19.245 2.645 ;
      RECT  18.925 2.645 19.25 2.65 ;
      RECT  18.925 2.65 19.255 2.655 ;
      RECT  18.925 2.655 19.26 2.66 ;
      RECT  18.93 2.66 19.265 2.665 ;
      RECT  18.935 2.665 19.27 2.67 ;
      RECT  18.94 2.67 19.275 2.675 ;
      RECT  18.945 2.675 19.28 2.68 ;
      RECT  18.95 2.68 19.285 2.685 ;
      RECT  18.955 2.685 19.29 2.69 ;
      RECT  18.96 2.69 19.295 2.695 ;
      RECT  18.965 2.695 19.3 2.7 ;
      RECT  18.97 2.7 19.305 2.705 ;
      RECT  18.975 2.705 19.31 2.71 ;
      RECT  18.98 2.71 19.315 2.715 ;
      RECT  18.985 2.715 19.32 2.72 ;
      RECT  18.99 2.72 19.325 2.725 ;
      RECT  18.995 2.725 19.33 2.73 ;
      RECT  19.0 2.73 19.335 2.735 ;
      RECT  19.005 2.735 19.34 2.74 ;
      RECT  19.01 2.74 19.345 2.745 ;
      RECT  19.015 2.745 19.35 2.75 ;
      RECT  19.02 2.75 19.355 2.755 ;
      RECT  19.025 2.755 19.36 2.76 ;
      RECT  19.03 2.76 19.365 2.765 ;
      RECT  19.035 2.765 19.37 2.77 ;
      RECT  19.04 2.77 19.375 2.775 ;
      RECT  19.045 2.775 19.38 2.78 ;
      RECT  19.05 2.78 19.385 2.785 ;
      RECT  19.055 2.785 19.39 2.79 ;
      RECT  19.06 2.79 19.395 2.795 ;
      RECT  19.065 2.795 19.4 2.8 ;
      RECT  19.07 2.8 19.405 2.805 ;
      RECT  19.075 2.805 19.41 2.81 ;
      RECT  19.08 2.81 19.415 2.815 ;
      RECT  19.085 2.815 19.42 2.82 ;
      RECT  19.09 2.82 19.425 2.825 ;
      RECT  19.095 2.825 19.43 2.83 ;
      RECT  19.1 2.83 19.435 2.835 ;
      RECT  19.105 2.835 19.44 2.84 ;
      RECT  19.11 2.84 19.445 2.845 ;
      RECT  19.115 2.845 19.45 2.85 ;
      RECT  19.12 2.85 19.455 2.855 ;
      RECT  19.125 2.855 19.46 2.86 ;
      RECT  19.13 2.86 19.465 2.865 ;
      RECT  19.135 2.865 19.47 2.87 ;
      RECT  19.14 2.87 19.475 2.875 ;
      RECT  19.145 2.875 19.48 2.88 ;
      RECT  19.15 2.88 19.485 2.885 ;
      RECT  19.155 2.885 19.49 2.89 ;
      RECT  19.16 2.89 19.495 2.895 ;
      RECT  19.165 2.895 19.5 2.9 ;
      RECT  19.17 2.9 19.505 2.905 ;
      RECT  19.175 2.905 19.51 2.91 ;
      RECT  19.18 2.91 19.515 2.915 ;
      RECT  19.185 2.915 19.52 2.92 ;
      RECT  19.19 2.92 19.525 2.925 ;
      RECT  19.195 2.925 19.53 2.93 ;
      RECT  19.2 2.93 19.535 2.935 ;
      RECT  19.205 2.935 19.54 2.94 ;
      RECT  19.21 2.94 19.545 2.945 ;
      RECT  19.215 2.945 19.55 2.95 ;
      RECT  19.22 2.95 19.555 2.955 ;
      RECT  19.225 2.955 19.56 2.96 ;
      RECT  19.23 2.96 19.565 2.965 ;
      RECT  19.235 2.965 19.57 2.97 ;
      RECT  19.24 2.97 19.575 2.975 ;
      RECT  19.245 2.975 19.58 2.98 ;
      RECT  19.25 2.98 19.585 2.985 ;
      RECT  19.255 2.985 19.59 2.99 ;
      RECT  19.26 2.99 19.595 2.995 ;
      RECT  19.265 2.995 19.6 3.0 ;
      RECT  19.27 3.0 19.605 3.005 ;
      RECT  19.275 3.005 19.61 3.01 ;
      RECT  19.28 3.01 19.615 3.015 ;
      RECT  19.285 3.015 19.62 3.02 ;
      RECT  19.29 3.02 19.625 3.025 ;
      RECT  19.295 3.025 19.63 3.03 ;
      RECT  19.3 3.03 19.635 3.035 ;
      RECT  19.305 3.035 19.64 3.04 ;
      RECT  19.31 3.04 19.645 3.045 ;
      RECT  19.315 3.045 19.65 3.05 ;
      RECT  19.32 3.05 19.655 3.055 ;
      RECT  19.325 3.055 19.66 3.06 ;
      RECT  19.33 3.06 19.665 3.065 ;
      RECT  19.335 3.065 19.67 3.07 ;
      RECT  19.34 3.07 19.675 3.075 ;
      RECT  19.345 3.075 19.68 3.08 ;
      RECT  19.35 3.08 19.685 3.085 ;
      RECT  19.355 3.085 19.69 3.09 ;
      RECT  19.36 3.09 19.695 3.095 ;
      RECT  19.365 3.095 19.7 3.1 ;
      RECT  19.37 3.1 19.705 3.105 ;
      RECT  19.375 3.105 19.71 3.11 ;
      RECT  19.38 3.11 19.715 3.115 ;
      RECT  19.385 3.115 19.715 3.12 ;
      RECT  19.39 3.12 19.715 3.125 ;
      RECT  19.395 3.125 19.715 3.13 ;
      RECT  19.4 3.13 19.715 3.135 ;
      RECT  19.405 3.135 19.715 3.14 ;
      RECT  19.41 3.14 19.715 3.145 ;
      RECT  19.415 3.145 19.715 3.15 ;
      RECT  19.42 3.15 19.715 3.155 ;
      RECT  19.425 3.155 19.715 3.16 ;
      RECT  19.43 3.16 19.715 3.165 ;
      RECT  19.435 3.165 19.715 3.17 ;
      RECT  19.44 3.17 19.715 3.175 ;
      RECT  19.445 3.175 19.715 3.18 ;
      RECT  19.45 3.18 19.715 3.185 ;
      RECT  19.455 3.185 19.715 3.19 ;
      RECT  19.46 3.19 19.715 3.195 ;
      RECT  19.465 3.195 19.715 3.2 ;
      RECT  19.47 3.2 19.715 3.205 ;
      RECT  19.475 3.205 19.715 3.21 ;
      RECT  19.48 3.21 19.715 3.215 ;
      RECT  19.485 3.215 19.715 3.81 ;
      RECT  16.94 3.7 18.475 3.81 ;
      RECT  16.94 3.81 19.715 3.93 ;
      RECT  18.245 3.93 19.715 4.04 ;
      RECT  16.94 3.93 17.17 4.155 ;
      RECT  13.62 4.155 17.17 4.385 ;
      RECT  4.015 1.61 4.245 1.89 ;
      RECT  4.015 1.89 4.595 2.12 ;
      RECT  4.365 2.12 4.595 2.405 ;
      RECT  4.365 2.405 5.21 2.635 ;
      RECT  4.365 2.635 4.595 3.245 ;
      RECT  3.96 3.245 4.595 3.475 ;
      RECT  5.485 3.81 8.515 4.04 ;
      RECT  5.485 4.04 5.715 4.365 ;
      RECT  8.285 4.04 8.515 4.465 ;
      RECT  4.66 4.365 5.715 4.595 ;
      RECT  8.285 4.465 11.02 4.695 ;
      RECT  9.14 4.005 13.26 4.235 ;
      RECT  17.4 4.16 18.035 4.39 ;
      RECT  17.805 4.39 18.035 4.54 ;
      RECT  17.805 4.54 19.155 4.77 ;
      RECT  18.925 4.77 19.155 5.0 ;
      RECT  18.925 5.0 20.89 5.23 ;
      RECT  0.18 4.365 1.74 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  19.64 4.365 22.22 4.595 ;
      RECT  11.645 4.62 17.475 4.85 ;
      RECT  11.645 4.85 11.875 5.0 ;
      RECT  17.245 4.85 17.475 5.0 ;
      RECT  9.35 5.0 11.875 5.155 ;
      RECT  17.245 5.0 18.65 5.23 ;
      RECT  9.35 5.155 11.87 5.23 ;
      RECT  3.75 5.0 7.45 5.23 ;
      LAYER METAL2 ;
      RECT  1.315 0.98 21.235 1.26 ;
      LAYER VIA12 ;
      RECT  1.375 0.99 1.635 1.25 ;
      RECT  9.95 0.99 10.21 1.25 ;
      RECT  20.915 0.99 21.175 1.25 ;
  END
END MDN_FSDNRBSBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNRBSBQ_2
#      Description : D-Flip Flop w/scan, neg-edge triggered, lo-async-clear/set, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNRBSBQ_2
  CLASS CORE ;
  FOREIGN MDN_FSDNRBSBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 24.64 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 8.54 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  22.58 1.565 24.46 1.795 ;
      RECT  23.405 1.795 23.635 3.245 ;
      RECT  22.575 3.245 24.46 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.325 2.125 16.38 2.355 ;
      RECT  13.325 2.355 13.555 2.38 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  13.25 2.38 13.555 2.405 ;
      RECT  12.71 2.405 13.555 2.635 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  21.7 4.365 21.98 5.0 ;
      RECT  21.67 5.0 22.01 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.81 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  20.72 5.46 21.395 5.74 ;
      RECT  16.63 5.09 16.97 5.46 ;
      RECT  16.24 5.46 17.36 5.74 ;
      RECT  12.15 5.09 12.49 5.46 ;
      RECT  11.76 5.46 15.12 5.74 ;
      RECT  14.39 5.09 14.73 5.46 ;
      RECT  6.2 4.365 7.955 4.595 ;
      RECT  7.725 4.595 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 24.64 5.74 ;
      LAYER VIA12 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  24.23 5.47 24.49 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 -0.14 24.81 0.14 ;
      RECT  23.405 0.14 23.635 0.73 ;
      RECT  21.84 -0.14 22.96 0.14 ;
      RECT  22.285 0.14 22.515 1.005 ;
      RECT  21.88 1.005 22.515 1.235 ;
      RECT  13.27 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 1.005 ;
      RECT  12.92 1.005 16.2 1.235 ;
      RECT  5.04 -0.14 6.16 0.14 ;
      RECT  5.43 0.14 5.77 0.465 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 24.64 0.14 ;
      LAYER VIA12 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  22.55 -0.13 22.81 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 10.81 0.445 ;
      RECT  6.045 0.445 10.81 0.675 ;
      RECT  6.045 0.675 6.275 0.695 ;
      RECT  3.805 0.445 5.155 0.675 ;
      RECT  4.925 0.675 5.155 0.695 ;
      RECT  3.805 0.675 4.035 1.005 ;
      RECT  4.925 0.695 6.275 0.925 ;
      RECT  2.63 0.37 2.97 0.6 ;
      RECT  2.63 0.6 2.86 1.005 ;
      RECT  1.565 1.005 4.035 1.235 ;
      RECT  1.565 1.235 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  12.205 0.37 14.19 0.6 ;
      RECT  12.205 0.6 12.435 1.465 ;
      RECT  9.965 1.465 12.435 1.695 ;
      RECT  9.965 1.695 10.195 3.53 ;
      RECT  14.95 0.37 22.01 0.6 ;
      RECT  23.91 0.37 24.25 0.6 ;
      RECT  23.91 0.6 24.14 1.005 ;
      RECT  22.79 0.37 23.13 0.6 ;
      RECT  22.9 0.6 23.13 1.005 ;
      RECT  22.9 1.005 24.14 1.235 ;
      RECT  17.51 0.83 21.395 1.06 ;
      RECT  17.51 1.06 17.74 1.565 ;
      RECT  21.165 1.06 21.395 2.405 ;
      RECT  16.685 1.565 17.74 1.795 ;
      RECT  16.685 1.795 16.915 3.245 ;
      RECT  20.55 2.405 23.005 2.635 ;
      RECT  15.86 3.245 17.74 3.475 ;
      RECT  6.605 1.005 8.78 1.155 ;
      RECT  4.66 1.155 8.78 1.235 ;
      RECT  4.66 1.235 6.835 1.385 ;
      RECT  10.68 1.005 11.72 1.235 ;
      RECT  18.1 1.29 20.68 1.52 ;
      RECT  3.96 1.565 4.3 1.62 ;
      RECT  3.96 1.62 4.595 1.85 ;
      RECT  4.365 1.85 4.595 2.41 ;
      RECT  4.365 2.41 5.21 2.64 ;
      RECT  4.365 2.64 4.595 3.245 ;
      RECT  3.96 3.245 4.595 3.475 ;
      RECT  7.67 1.565 9.48 1.795 ;
      RECT  6.2 1.615 7.24 1.845 ;
      RECT  18.87 1.75 19.21 1.98 ;
      RECT  18.925 1.98 19.155 2.405 ;
      RECT  17.19 2.405 19.155 2.635 ;
      RECT  18.925 2.635 19.155 3.48 ;
      RECT  19.485 1.75 19.98 1.98 ;
      RECT  19.485 1.98 19.715 3.71 ;
      RECT  12.765 1.565 13.96 1.795 ;
      RECT  12.765 1.795 12.995 1.94 ;
      RECT  11.645 1.94 12.995 2.17 ;
      RECT  11.645 2.17 11.875 3.03 ;
      RECT  11.645 3.03 14.675 3.26 ;
      RECT  14.445 3.26 14.675 3.71 ;
      RECT  14.445 3.71 19.715 3.94 ;
      RECT  4.925 3.245 8.91 3.475 ;
      RECT  4.925 3.475 5.155 3.805 ;
      RECT  8.68 3.475 8.91 4.48 ;
      RECT  4.66 3.805 5.155 4.035 ;
      RECT  8.68 4.48 11.02 4.71 ;
      RECT  20.045 3.245 22.22 3.475 ;
      RECT  20.045 3.475 20.275 4.365 ;
      RECT  19.64 4.365 20.275 4.595 ;
      RECT  10.525 2.35 10.755 3.49 ;
      RECT  10.525 3.49 14.115 3.72 ;
      RECT  13.885 3.72 14.115 4.17 ;
      RECT  13.885 4.17 19.155 4.4 ;
      RECT  18.925 4.4 19.155 5.0 ;
      RECT  18.925 5.0 19.77 5.23 ;
      RECT  9.14 3.95 13.26 4.18 ;
      RECT  11.645 4.63 18.5 4.86 ;
      RECT  11.645 4.86 11.875 5.0 ;
      RECT  18.27 4.86 18.5 5.0 ;
      RECT  5.485 3.805 8.42 4.035 ;
      RECT  5.485 4.035 5.715 4.365 ;
      RECT  8.19 4.035 8.42 5.0 ;
      RECT  2.42 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  2.42 3.245 2.915 3.475 ;
      RECT  2.685 3.475 2.915 4.365 ;
      RECT  2.685 4.365 5.715 4.595 ;
      RECT  8.19 5.0 11.875 5.23 ;
      RECT  18.27 5.0 18.65 5.23 ;
      RECT  3.75 5.0 7.45 5.23 ;
  END
END MDN_FSDNRBSBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNRBSBQ_4
#      Description : D-Flip Flop w/scan, neg-edge triggered, lo-async-clear/set, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNRBSBQ_4
  CLASS CORE ;
  FOREIGN MDN_FSDNRBSBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 26.88 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 8.54 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  22.58 1.565 26.7 1.795 ;
      RECT  24.525 1.795 24.755 3.245 ;
      RECT  22.57 3.245 26.7 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.325 2.125 16.38 2.355 ;
      RECT  13.325 2.355 13.555 2.38 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  13.25 2.38 13.555 2.405 ;
      RECT  12.71 2.405 13.555 2.635 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  21.7 4.365 21.98 5.0 ;
      RECT  21.67 5.0 22.01 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.645 5.46 27.05 5.74 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.08 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  20.72 5.46 21.395 5.74 ;
      RECT  14.39 5.135 14.73 5.46 ;
      RECT  14.0 5.46 17.36 5.74 ;
      RECT  16.63 5.135 16.97 5.46 ;
      RECT  12.15 5.135 12.49 5.46 ;
      RECT  11.76 5.46 12.88 5.74 ;
      RECT  6.2 4.48 7.955 4.71 ;
      RECT  7.725 4.71 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 26.88 5.74 ;
      LAYER VIA12 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 -0.14 27.05 0.14 ;
      RECT  25.645 0.14 25.875 0.7 ;
      RECT  22.96 -0.14 24.08 0.14 ;
      RECT  23.405 0.14 23.635 1.005 ;
      RECT  21.88 1.005 23.635 1.235 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 1.005 ;
      RECT  12.92 1.005 16.2 1.235 ;
      RECT  5.04 -0.14 6.16 0.14 ;
      RECT  5.43 0.14 5.77 0.465 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.66 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 26.88 0.14 ;
      LAYER VIA12 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  23.11 -0.13 23.37 0.13 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  13.83 0.37 14.17 0.445 ;
      RECT  12.205 0.445 14.17 0.675 ;
      RECT  12.205 0.675 12.435 1.48 ;
      RECT  9.965 1.48 12.435 1.71 ;
      RECT  9.965 1.71 10.195 3.53 ;
      RECT  9.965 0.37 10.81 0.6 ;
      RECT  9.965 0.6 10.195 0.74 ;
      RECT  3.805 0.74 10.195 0.97 ;
      RECT  3.805 0.97 4.035 1.005 ;
      RECT  2.63 0.37 2.97 0.6 ;
      RECT  2.63 0.6 2.86 1.005 ;
      RECT  1.565 1.005 4.035 1.235 ;
      RECT  1.565 1.235 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  14.95 0.37 22.01 0.6 ;
      RECT  17.51 0.83 21.395 1.06 ;
      RECT  17.51 1.06 17.74 1.565 ;
      RECT  21.165 1.06 21.395 2.125 ;
      RECT  16.685 1.565 17.74 1.795 ;
      RECT  16.685 1.795 16.915 3.245 ;
      RECT  20.605 2.125 24.195 2.355 ;
      RECT  20.605 2.355 20.835 2.69 ;
      RECT  22.845 2.355 23.075 2.69 ;
      RECT  23.965 2.355 24.195 2.69 ;
      RECT  15.86 3.245 17.74 3.475 ;
      RECT  10.68 1.005 11.72 1.235 ;
      RECT  4.66 1.2 8.78 1.43 ;
      RECT  18.1 1.29 20.68 1.52 ;
      RECT  3.96 1.655 4.595 1.885 ;
      RECT  4.365 1.885 4.595 2.405 ;
      RECT  4.365 2.405 5.215 2.635 ;
      RECT  4.365 2.635 4.595 3.245 ;
      RECT  3.91 3.245 4.595 3.475 ;
      RECT  6.2 1.66 7.24 1.89 ;
      RECT  7.67 1.66 9.48 1.89 ;
      RECT  18.365 1.75 19.16 1.98 ;
      RECT  18.365 1.98 18.595 2.405 ;
      RECT  17.19 2.405 18.595 2.635 ;
      RECT  18.365 2.635 18.595 3.245 ;
      RECT  18.365 3.245 19.16 3.475 ;
      RECT  19.485 1.75 19.98 1.98 ;
      RECT  19.485 1.98 19.715 3.755 ;
      RECT  12.765 1.565 13.96 1.795 ;
      RECT  12.765 1.795 12.995 1.94 ;
      RECT  11.645 1.94 12.995 2.17 ;
      RECT  11.645 2.17 11.875 3.03 ;
      RECT  11.645 3.03 14.675 3.26 ;
      RECT  14.445 3.26 14.675 3.755 ;
      RECT  14.445 3.755 19.715 3.985 ;
      RECT  25.085 2.125 26.435 2.355 ;
      RECT  25.085 2.355 25.315 2.685 ;
      RECT  26.205 2.355 26.435 2.685 ;
      RECT  4.925 3.245 8.875 3.475 ;
      RECT  4.925 3.475 5.155 3.805 ;
      RECT  8.645 3.475 8.875 4.48 ;
      RECT  4.66 3.805 5.155 4.035 ;
      RECT  8.645 4.48 11.02 4.71 ;
      RECT  20.045 3.245 22.22 3.475 ;
      RECT  20.045 3.475 20.275 4.365 ;
      RECT  19.635 4.365 20.275 4.595 ;
      RECT  10.525 2.35 10.755 3.56 ;
      RECT  10.525 3.56 14.115 3.79 ;
      RECT  13.885 3.79 14.115 4.215 ;
      RECT  13.885 4.215 19.155 4.445 ;
      RECT  18.925 4.445 19.155 5.0 ;
      RECT  18.925 5.0 19.77 5.23 ;
      RECT  9.14 4.02 13.26 4.25 ;
      RECT  11.645 4.675 18.52 4.905 ;
      RECT  11.645 4.905 11.875 5.0 ;
      RECT  18.29 4.905 18.52 5.0 ;
      RECT  5.485 3.805 8.415 4.035 ;
      RECT  5.485 4.035 5.715 4.365 ;
      RECT  8.185 4.035 8.415 5.0 ;
      RECT  2.42 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  2.42 3.245 2.915 3.475 ;
      RECT  2.685 3.475 2.915 4.365 ;
      RECT  2.685 4.365 5.715 4.595 ;
      RECT  8.185 5.0 11.875 5.23 ;
      RECT  18.29 5.0 18.65 5.23 ;
      RECT  3.75 5.0 7.45 5.23 ;
      RECT  23.91 5.0 25.37 5.23 ;
  END
END MDN_FSDNRBSBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNSBQ_1
#      Description : D-Flip Flop w/scan, neg-edge triggered, lo-async-/set, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNSBQ_1
  CLASS CORE ;
  FOREIGN MDN_FSDNSBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 1.565 9.66 2.355 ;
      RECT  9.405 2.355 9.635 2.69 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.54 0.6 1.82 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.485 1.565 19.98 1.795 ;
      RECT  19.485 1.795 19.715 3.245 ;
      RECT  19.485 3.245 19.98 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.98 2.125 17.5 2.355 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.63 5.135 16.97 5.46 ;
      RECT  16.24 5.46 17.36 5.74 ;
      RECT  14.39 5.135 14.73 5.46 ;
      RECT  14.0 5.46 15.12 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 11.37 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.19 5.135 3.53 5.46 ;
      RECT  2.8 5.46 3.92 5.74 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  15.12 -0.14 15.85 0.14 ;
      RECT  15.565 0.14 15.795 1.005 ;
      RECT  15.16 1.005 17.74 1.235 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.685 -0.14 3.36 0.14 ;
      RECT  2.685 0.14 2.915 1.005 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 10.81 0.445 ;
      RECT  10.47 0.445 13.05 0.675 ;
      RECT  12.71 0.37 13.05 0.445 ;
      RECT  10.47 0.675 10.7 1.005 ;
      RECT  7.11 0.37 7.45 0.445 ;
      RECT  7.11 0.445 9.37 0.675 ;
      RECT  9.14 0.675 9.37 1.005 ;
      RECT  9.14 1.005 10.7 1.235 ;
      RECT  9.965 1.235 10.195 3.05 ;
      RECT  9.14 3.05 10.195 3.28 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  19.43 0.37 19.77 0.6 ;
      RECT  19.43 0.6 19.66 1.005 ;
      RECT  16.07 0.37 16.41 0.445 ;
      RECT  16.07 0.445 18.29 0.675 ;
      RECT  18.06 0.675 18.29 1.005 ;
      RECT  18.06 1.005 19.66 1.235 ;
      RECT  18.365 1.235 18.595 3.245 ;
      RECT  18.1 3.245 18.595 3.475 ;
      RECT  11.38 1.005 14.6 1.01 ;
      RECT  11.38 1.01 14.605 1.015 ;
      RECT  11.38 1.015 14.61 1.02 ;
      RECT  11.38 1.02 14.615 1.025 ;
      RECT  11.38 1.025 14.62 1.03 ;
      RECT  11.38 1.03 14.625 1.035 ;
      RECT  11.38 1.035 14.63 1.04 ;
      RECT  11.38 1.04 14.635 1.045 ;
      RECT  11.38 1.045 14.64 1.05 ;
      RECT  11.38 1.05 14.645 1.055 ;
      RECT  11.38 1.055 14.65 1.06 ;
      RECT  11.38 1.06 14.655 1.065 ;
      RECT  11.38 1.065 14.66 1.07 ;
      RECT  11.38 1.07 14.665 1.075 ;
      RECT  11.38 1.075 14.67 1.08 ;
      RECT  11.38 1.08 14.675 1.085 ;
      RECT  11.38 1.085 14.68 1.09 ;
      RECT  11.38 1.09 14.685 1.095 ;
      RECT  11.38 1.095 14.69 1.1 ;
      RECT  11.38 1.1 14.695 1.105 ;
      RECT  11.38 1.105 14.7 1.11 ;
      RECT  11.38 1.11 14.705 1.115 ;
      RECT  11.38 1.115 14.71 1.12 ;
      RECT  11.38 1.12 14.715 1.125 ;
      RECT  11.38 1.125 14.72 1.13 ;
      RECT  11.38 1.13 14.725 1.135 ;
      RECT  11.38 1.135 14.73 1.14 ;
      RECT  11.38 1.14 14.735 1.145 ;
      RECT  11.38 1.145 14.74 1.15 ;
      RECT  11.38 1.15 14.745 1.155 ;
      RECT  11.38 1.155 14.75 1.16 ;
      RECT  11.38 1.16 14.755 1.165 ;
      RECT  11.38 1.165 14.76 1.17 ;
      RECT  11.38 1.17 14.765 1.175 ;
      RECT  11.38 1.175 14.77 1.18 ;
      RECT  11.38 1.18 14.775 1.185 ;
      RECT  11.38 1.185 14.78 1.19 ;
      RECT  11.38 1.19 14.785 1.195 ;
      RECT  11.38 1.195 14.79 1.2 ;
      RECT  11.38 1.2 14.795 1.205 ;
      RECT  11.38 1.205 14.8 1.21 ;
      RECT  11.38 1.21 14.805 1.215 ;
      RECT  11.38 1.215 14.81 1.22 ;
      RECT  11.38 1.22 14.815 1.225 ;
      RECT  11.38 1.225 14.82 1.23 ;
      RECT  11.38 1.23 14.825 1.235 ;
      RECT  14.495 1.235 14.83 1.24 ;
      RECT  14.5 1.24 14.835 1.245 ;
      RECT  14.505 1.245 14.84 1.25 ;
      RECT  14.51 1.25 14.845 1.255 ;
      RECT  14.515 1.255 14.85 1.26 ;
      RECT  14.52 1.26 14.855 1.265 ;
      RECT  14.525 1.265 14.86 1.27 ;
      RECT  14.53 1.27 14.865 1.275 ;
      RECT  14.535 1.275 14.87 1.28 ;
      RECT  14.54 1.28 14.875 1.285 ;
      RECT  14.545 1.285 14.88 1.29 ;
      RECT  14.55 1.29 14.885 1.295 ;
      RECT  14.555 1.295 14.89 1.3 ;
      RECT  14.56 1.3 14.895 1.305 ;
      RECT  14.565 1.305 14.9 1.31 ;
      RECT  14.57 1.31 14.905 1.315 ;
      RECT  14.575 1.315 14.91 1.32 ;
      RECT  14.58 1.32 14.915 1.325 ;
      RECT  14.585 1.325 14.92 1.33 ;
      RECT  14.59 1.33 14.925 1.335 ;
      RECT  14.595 1.335 14.93 1.34 ;
      RECT  14.6 1.34 14.935 1.345 ;
      RECT  14.605 1.345 14.94 1.35 ;
      RECT  14.61 1.35 14.945 1.355 ;
      RECT  14.615 1.355 14.95 1.36 ;
      RECT  14.62 1.36 14.955 1.365 ;
      RECT  14.625 1.365 14.96 1.37 ;
      RECT  14.63 1.37 14.965 1.375 ;
      RECT  14.635 1.375 14.97 1.38 ;
      RECT  14.64 1.38 14.975 1.385 ;
      RECT  14.645 1.385 14.98 1.39 ;
      RECT  14.65 1.39 14.985 1.395 ;
      RECT  14.655 1.395 14.99 1.4 ;
      RECT  14.66 1.4 14.995 1.405 ;
      RECT  14.665 1.405 15.0 1.41 ;
      RECT  14.67 1.41 15.005 1.415 ;
      RECT  14.675 1.415 15.01 1.42 ;
      RECT  14.68 1.42 15.015 1.425 ;
      RECT  14.685 1.425 15.02 1.43 ;
      RECT  14.69 1.43 15.025 1.435 ;
      RECT  14.695 1.435 15.03 1.44 ;
      RECT  14.7 1.44 15.035 1.445 ;
      RECT  14.705 1.445 15.04 1.45 ;
      RECT  14.71 1.45 15.045 1.455 ;
      RECT  14.715 1.455 15.05 1.46 ;
      RECT  14.72 1.46 15.055 1.465 ;
      RECT  14.725 1.465 15.06 1.47 ;
      RECT  14.73 1.47 15.065 1.475 ;
      RECT  14.735 1.475 15.07 1.48 ;
      RECT  14.74 1.48 15.075 1.485 ;
      RECT  14.745 1.485 15.08 1.49 ;
      RECT  14.75 1.49 15.085 1.495 ;
      RECT  14.755 1.495 15.09 1.5 ;
      RECT  14.76 1.5 15.095 1.505 ;
      RECT  14.765 1.505 15.1 1.51 ;
      RECT  14.77 1.51 15.105 1.515 ;
      RECT  14.775 1.515 15.11 1.52 ;
      RECT  14.78 1.52 15.115 1.525 ;
      RECT  14.785 1.525 15.12 1.53 ;
      RECT  14.79 1.53 15.125 1.535 ;
      RECT  14.795 1.535 15.13 1.54 ;
      RECT  14.8 1.54 15.135 1.545 ;
      RECT  14.805 1.545 15.14 1.55 ;
      RECT  14.81 1.55 15.145 1.555 ;
      RECT  14.815 1.555 15.15 1.56 ;
      RECT  14.82 1.56 15.155 1.565 ;
      RECT  14.825 1.565 16.2 1.57 ;
      RECT  14.83 1.57 16.2 1.575 ;
      RECT  14.835 1.575 16.2 1.58 ;
      RECT  14.84 1.58 16.2 1.585 ;
      RECT  14.845 1.585 16.2 1.59 ;
      RECT  14.85 1.59 16.2 1.595 ;
      RECT  14.855 1.595 16.2 1.6 ;
      RECT  14.86 1.6 16.2 1.605 ;
      RECT  14.865 1.605 16.2 1.61 ;
      RECT  14.87 1.61 16.2 1.615 ;
      RECT  14.875 1.615 16.2 1.62 ;
      RECT  14.88 1.62 16.2 1.625 ;
      RECT  14.885 1.625 16.2 1.63 ;
      RECT  14.89 1.63 16.2 1.635 ;
      RECT  14.895 1.635 16.2 1.64 ;
      RECT  14.9 1.64 16.2 1.645 ;
      RECT  14.905 1.645 16.2 1.65 ;
      RECT  14.91 1.65 16.2 1.655 ;
      RECT  14.915 1.655 16.2 1.66 ;
      RECT  14.92 1.66 16.2 1.665 ;
      RECT  14.925 1.665 16.2 1.67 ;
      RECT  14.93 1.67 16.2 1.675 ;
      RECT  14.935 1.675 16.2 1.68 ;
      RECT  14.94 1.68 16.2 1.685 ;
      RECT  14.945 1.685 16.2 1.69 ;
      RECT  14.95 1.69 16.2 1.695 ;
      RECT  14.955 1.695 16.2 1.7 ;
      RECT  14.96 1.7 16.2 1.705 ;
      RECT  14.965 1.705 16.2 1.71 ;
      RECT  14.97 1.71 16.2 1.715 ;
      RECT  14.975 1.715 16.2 1.72 ;
      RECT  14.98 1.72 16.2 1.725 ;
      RECT  14.985 1.725 16.2 1.73 ;
      RECT  14.99 1.73 16.2 1.735 ;
      RECT  14.995 1.735 16.2 1.74 ;
      RECT  15.0 1.74 16.2 1.745 ;
      RECT  15.005 1.745 16.2 1.75 ;
      RECT  15.01 1.75 16.2 1.755 ;
      RECT  15.015 1.755 16.2 1.76 ;
      RECT  15.02 1.76 16.2 1.765 ;
      RECT  15.025 1.765 16.2 1.77 ;
      RECT  15.03 1.77 16.2 1.775 ;
      RECT  15.035 1.775 16.2 1.78 ;
      RECT  15.04 1.78 16.2 1.785 ;
      RECT  15.045 1.785 16.2 1.79 ;
      RECT  15.05 1.79 16.2 1.795 ;
      RECT  3.24 1.005 8.78 1.235 ;
      RECT  3.24 1.235 3.48 1.565 ;
      RECT  1.715 1.565 3.48 1.795 ;
      RECT  4.365 1.565 5.0 1.795 ;
      RECT  4.365 1.795 4.595 3.75 ;
      RECT  0.49 3.75 5.0 3.98 ;
      RECT  0.49 3.98 0.72 5.0 ;
      RECT  0.38 5.0 0.72 5.23 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  10.68 1.565 11.315 1.795 ;
      RECT  11.085 1.795 11.315 2.425 ;
      RECT  11.085 2.425 11.93 2.655 ;
      RECT  11.085 2.655 11.315 3.245 ;
      RECT  10.68 3.245 11.315 3.475 ;
      RECT  12.92 1.75 14.675 1.98 ;
      RECT  14.445 1.98 14.675 3.755 ;
      RECT  13.26 3.755 15.5 3.76 ;
      RECT  13.255 3.76 15.5 3.765 ;
      RECT  13.25 3.765 15.5 3.77 ;
      RECT  13.245 3.77 15.5 3.775 ;
      RECT  13.24 3.775 15.5 3.78 ;
      RECT  13.235 3.78 15.5 3.785 ;
      RECT  13.23 3.785 15.5 3.79 ;
      RECT  13.225 3.79 15.5 3.795 ;
      RECT  13.22 3.795 15.5 3.8 ;
      RECT  13.215 3.8 15.5 3.805 ;
      RECT  13.21 3.805 15.5 3.81 ;
      RECT  13.205 3.81 15.5 3.815 ;
      RECT  13.2 3.815 15.5 3.82 ;
      RECT  13.195 3.82 15.5 3.825 ;
      RECT  13.19 3.825 15.5 3.83 ;
      RECT  13.185 3.83 15.5 3.835 ;
      RECT  13.18 3.835 15.5 3.84 ;
      RECT  13.175 3.84 15.5 3.845 ;
      RECT  13.17 3.845 15.5 3.85 ;
      RECT  13.165 3.85 15.5 3.855 ;
      RECT  13.16 3.855 15.5 3.86 ;
      RECT  13.155 3.86 15.5 3.865 ;
      RECT  13.15 3.865 15.5 3.87 ;
      RECT  13.145 3.87 15.5 3.875 ;
      RECT  13.14 3.875 15.5 3.88 ;
      RECT  13.135 3.88 15.5 3.885 ;
      RECT  13.13 3.885 15.5 3.89 ;
      RECT  13.125 3.89 15.5 3.895 ;
      RECT  13.12 3.895 15.5 3.9 ;
      RECT  13.115 3.9 15.5 3.905 ;
      RECT  13.11 3.905 15.5 3.91 ;
      RECT  13.105 3.91 15.5 3.915 ;
      RECT  13.1 3.915 15.5 3.92 ;
      RECT  13.095 3.92 15.5 3.925 ;
      RECT  13.09 3.925 15.5 3.93 ;
      RECT  13.085 3.93 15.5 3.935 ;
      RECT  13.08 3.935 15.5 3.94 ;
      RECT  13.075 3.94 15.5 3.945 ;
      RECT  13.07 3.945 15.5 3.95 ;
      RECT  13.065 3.95 15.5 3.955 ;
      RECT  13.06 3.955 15.5 3.96 ;
      RECT  13.055 3.96 15.5 3.965 ;
      RECT  13.05 3.965 15.5 3.97 ;
      RECT  13.045 3.97 15.5 3.975 ;
      RECT  13.04 3.975 15.5 3.98 ;
      RECT  13.035 3.98 15.5 3.985 ;
      RECT  13.03 3.985 13.355 3.99 ;
      RECT  13.025 3.99 13.35 3.995 ;
      RECT  13.02 3.995 13.345 4.0 ;
      RECT  13.015 4.0 13.34 4.005 ;
      RECT  13.01 4.005 13.335 4.01 ;
      RECT  13.005 4.01 13.33 4.015 ;
      RECT  13.0 4.015 13.325 4.02 ;
      RECT  12.205 4.02 13.32 4.025 ;
      RECT  12.205 4.025 13.315 4.03 ;
      RECT  12.205 4.03 13.31 4.035 ;
      RECT  12.205 4.035 13.305 4.04 ;
      RECT  12.205 4.04 13.3 4.045 ;
      RECT  12.205 4.045 13.295 4.05 ;
      RECT  12.205 4.05 13.29 4.055 ;
      RECT  12.205 4.055 13.285 4.06 ;
      RECT  12.205 4.06 13.28 4.065 ;
      RECT  12.205 4.065 13.275 4.07 ;
      RECT  12.205 4.07 13.27 4.075 ;
      RECT  12.205 4.075 13.265 4.08 ;
      RECT  12.205 4.08 13.26 4.085 ;
      RECT  12.205 4.085 13.255 4.09 ;
      RECT  12.205 4.09 13.25 4.095 ;
      RECT  12.205 4.095 13.245 4.1 ;
      RECT  12.205 4.1 13.24 4.105 ;
      RECT  12.205 4.105 13.235 4.11 ;
      RECT  12.205 4.11 13.23 4.115 ;
      RECT  12.205 4.115 13.225 4.12 ;
      RECT  12.205 4.12 13.22 4.125 ;
      RECT  12.205 4.125 13.215 4.13 ;
      RECT  12.205 4.13 13.21 4.135 ;
      RECT  12.205 4.135 13.205 4.14 ;
      RECT  12.205 4.14 13.2 4.145 ;
      RECT  12.205 4.145 13.195 4.15 ;
      RECT  12.205 4.15 13.19 4.155 ;
      RECT  12.205 4.155 13.185 4.16 ;
      RECT  12.205 4.16 13.18 4.165 ;
      RECT  12.205 4.165 13.175 4.17 ;
      RECT  12.205 4.17 13.17 4.175 ;
      RECT  12.205 4.175 13.165 4.18 ;
      RECT  12.205 4.18 13.16 4.185 ;
      RECT  12.205 4.185 13.155 4.19 ;
      RECT  12.205 4.19 13.15 4.195 ;
      RECT  12.205 4.195 13.145 4.2 ;
      RECT  12.205 4.2 13.14 4.205 ;
      RECT  8.955 4.205 13.135 4.21 ;
      RECT  8.955 4.21 13.13 4.215 ;
      RECT  8.955 4.215 13.125 4.22 ;
      RECT  8.955 4.22 13.12 4.225 ;
      RECT  8.955 4.225 13.115 4.23 ;
      RECT  8.955 4.23 13.11 4.235 ;
      RECT  8.955 4.235 13.105 4.24 ;
      RECT  8.955 4.24 13.1 4.245 ;
      RECT  8.955 4.245 13.095 4.25 ;
      RECT  8.955 4.25 12.435 4.435 ;
      RECT  8.955 4.435 9.185 4.54 ;
      RECT  7.725 4.54 9.185 4.77 ;
      RECT  7.725 4.77 7.955 5.0 ;
      RECT  5.99 5.0 7.955 5.23 ;
      RECT  12.665 2.39 14.01 2.62 ;
      RECT  12.665 2.62 12.895 3.555 ;
      RECT  11.645 3.555 12.895 3.745 ;
      RECT  7.725 1.585 7.955 3.51 ;
      RECT  7.725 3.51 9.185 3.74 ;
      RECT  8.955 3.74 9.185 3.745 ;
      RECT  8.955 3.745 12.895 3.785 ;
      RECT  8.955 3.785 11.875 3.975 ;
      RECT  12.205 1.59 12.435 3.315 ;
      RECT  0.175 3.245 2.76 3.475 ;
      RECT  5.485 3.245 7.24 3.475 ;
      RECT  5.485 3.475 5.715 4.365 ;
      RECT  4.925 4.365 5.715 4.595 ;
      RECT  4.925 4.595 5.155 4.675 ;
      RECT  2.68 4.675 5.155 4.905 ;
      RECT  2.68 4.905 2.92 4.925 ;
      RECT  0.95 4.925 2.92 5.155 ;
      RECT  8.495 3.97 8.725 4.08 ;
      RECT  6.2 4.08 8.725 4.31 ;
      RECT  1.72 4.215 4.3 4.445 ;
      RECT  13.47 4.215 17.74 4.445 ;
      RECT  13.47 4.445 13.7 4.48 ;
      RECT  12.92 4.48 13.7 4.71 ;
      RECT  9.415 4.665 10.755 4.905 ;
      RECT  9.415 4.905 9.645 5.0 ;
      RECT  10.525 4.905 10.755 5.0 ;
      RECT  8.23 5.0 9.645 5.23 ;
      RECT  10.525 5.0 11.92 5.23 ;
      RECT  13.93 4.675 17.475 4.905 ;
      RECT  17.245 4.905 17.475 4.925 ;
      RECT  13.93 4.905 14.16 4.98 ;
      RECT  17.245 4.925 18.65 5.155 ;
      RECT  12.15 4.98 14.16 5.21 ;
      RECT  18.31 5.155 18.65 5.23 ;
  END
END MDN_FSDNSBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNSBQ_2
#      Description : D-Flip Flop w/scan, neg-edge triggered, lo-async-/set, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNSBQ_2
  CLASS CORE ;
  FOREIGN MDN_FSDNSBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 9.635 2.355 ;
      RECT  9.405 2.355 9.635 2.69 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.54 0.6 1.82 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.64 1.565 20.68 1.795 ;
      RECT  20.045 1.795 20.275 3.245 ;
      RECT  19.64 3.245 20.68 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.98 2.125 17.5 2.355 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.87 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  14.39 5.135 14.73 5.46 ;
      RECT  14.0 5.46 17.36 5.74 ;
      RECT  16.63 5.135 16.97 5.46 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 10.64 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.19 5.135 3.53 5.46 ;
      RECT  2.8 5.46 3.92 5.74 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  15.12 -0.14 16.24 0.14 ;
      RECT  15.565 0.14 15.795 1.005 ;
      RECT  15.16 1.005 17.74 1.235 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.685 -0.14 3.36 0.14 ;
      RECT  2.685 0.14 2.915 1.005 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 10.81 0.445 ;
      RECT  10.47 0.445 13.05 0.675 ;
      RECT  12.71 0.37 13.05 0.445 ;
      RECT  10.47 0.675 10.7 1.005 ;
      RECT  7.11 0.37 7.45 0.445 ;
      RECT  7.11 0.445 9.635 0.675 ;
      RECT  9.405 0.675 9.635 1.005 ;
      RECT  9.405 1.005 10.7 1.235 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  19.43 0.37 20.89 0.6 ;
      RECT  19.43 0.6 19.66 1.005 ;
      RECT  16.07 0.37 18.33 0.6 ;
      RECT  18.1 0.6 18.33 1.005 ;
      RECT  18.1 1.005 19.66 1.235 ;
      RECT  18.925 1.235 19.155 4.365 ;
      RECT  18.1 4.365 19.155 4.595 ;
      RECT  11.38 1.005 14.6 1.01 ;
      RECT  11.38 1.01 14.605 1.015 ;
      RECT  11.38 1.015 14.61 1.02 ;
      RECT  11.38 1.02 14.615 1.025 ;
      RECT  11.38 1.025 14.62 1.03 ;
      RECT  11.38 1.03 14.625 1.035 ;
      RECT  11.38 1.035 14.63 1.04 ;
      RECT  11.38 1.04 14.635 1.045 ;
      RECT  11.38 1.045 14.64 1.05 ;
      RECT  11.38 1.05 14.645 1.055 ;
      RECT  11.38 1.055 14.65 1.06 ;
      RECT  11.38 1.06 14.655 1.065 ;
      RECT  11.38 1.065 14.66 1.07 ;
      RECT  11.38 1.07 14.665 1.075 ;
      RECT  11.38 1.075 14.67 1.08 ;
      RECT  11.38 1.08 14.675 1.085 ;
      RECT  11.38 1.085 14.68 1.09 ;
      RECT  11.38 1.09 14.685 1.095 ;
      RECT  11.38 1.095 14.69 1.1 ;
      RECT  11.38 1.1 14.695 1.105 ;
      RECT  11.38 1.105 14.7 1.11 ;
      RECT  11.38 1.11 14.705 1.115 ;
      RECT  11.38 1.115 14.71 1.12 ;
      RECT  11.38 1.12 14.715 1.125 ;
      RECT  11.38 1.125 14.72 1.13 ;
      RECT  11.38 1.13 14.725 1.135 ;
      RECT  11.38 1.135 14.73 1.14 ;
      RECT  11.38 1.14 14.735 1.145 ;
      RECT  11.38 1.145 14.74 1.15 ;
      RECT  11.38 1.15 14.745 1.155 ;
      RECT  11.38 1.155 14.75 1.16 ;
      RECT  11.38 1.16 14.755 1.165 ;
      RECT  11.38 1.165 14.76 1.17 ;
      RECT  11.38 1.17 14.765 1.175 ;
      RECT  11.38 1.175 14.77 1.18 ;
      RECT  11.38 1.18 14.775 1.185 ;
      RECT  11.38 1.185 14.78 1.19 ;
      RECT  11.38 1.19 14.785 1.195 ;
      RECT  11.38 1.195 14.79 1.2 ;
      RECT  11.38 1.2 14.795 1.205 ;
      RECT  11.38 1.205 14.8 1.21 ;
      RECT  11.38 1.21 14.805 1.215 ;
      RECT  11.38 1.215 14.81 1.22 ;
      RECT  11.38 1.22 14.815 1.225 ;
      RECT  11.38 1.225 14.82 1.23 ;
      RECT  11.38 1.23 14.825 1.235 ;
      RECT  14.495 1.235 14.83 1.24 ;
      RECT  14.5 1.24 14.835 1.245 ;
      RECT  14.505 1.245 14.84 1.25 ;
      RECT  14.51 1.25 14.845 1.255 ;
      RECT  14.515 1.255 14.85 1.26 ;
      RECT  14.52 1.26 14.855 1.265 ;
      RECT  14.525 1.265 14.86 1.27 ;
      RECT  14.53 1.27 14.865 1.275 ;
      RECT  14.535 1.275 14.87 1.28 ;
      RECT  14.54 1.28 14.875 1.285 ;
      RECT  14.545 1.285 14.88 1.29 ;
      RECT  14.55 1.29 14.885 1.295 ;
      RECT  14.555 1.295 14.89 1.3 ;
      RECT  14.56 1.3 14.895 1.305 ;
      RECT  14.565 1.305 14.9 1.31 ;
      RECT  14.57 1.31 14.905 1.315 ;
      RECT  14.575 1.315 14.91 1.32 ;
      RECT  14.58 1.32 14.915 1.325 ;
      RECT  14.585 1.325 14.92 1.33 ;
      RECT  14.59 1.33 14.925 1.335 ;
      RECT  14.595 1.335 14.93 1.34 ;
      RECT  14.6 1.34 14.935 1.345 ;
      RECT  14.605 1.345 14.94 1.35 ;
      RECT  14.61 1.35 14.945 1.355 ;
      RECT  14.615 1.355 14.95 1.36 ;
      RECT  14.62 1.36 14.955 1.365 ;
      RECT  14.625 1.365 14.96 1.37 ;
      RECT  14.63 1.37 14.965 1.375 ;
      RECT  14.635 1.375 14.97 1.38 ;
      RECT  14.64 1.38 14.975 1.385 ;
      RECT  14.645 1.385 14.98 1.39 ;
      RECT  14.65 1.39 14.985 1.395 ;
      RECT  14.655 1.395 14.99 1.4 ;
      RECT  14.66 1.4 14.995 1.405 ;
      RECT  14.665 1.405 15.0 1.41 ;
      RECT  14.67 1.41 15.005 1.415 ;
      RECT  14.675 1.415 15.01 1.42 ;
      RECT  14.68 1.42 15.015 1.425 ;
      RECT  14.685 1.425 15.02 1.43 ;
      RECT  14.69 1.43 15.025 1.435 ;
      RECT  14.695 1.435 15.03 1.44 ;
      RECT  14.7 1.44 15.035 1.445 ;
      RECT  14.705 1.445 15.04 1.45 ;
      RECT  14.71 1.45 15.045 1.455 ;
      RECT  14.715 1.455 15.05 1.46 ;
      RECT  14.72 1.46 15.055 1.465 ;
      RECT  14.725 1.465 15.06 1.47 ;
      RECT  14.73 1.47 15.065 1.475 ;
      RECT  14.735 1.475 15.07 1.48 ;
      RECT  14.74 1.48 15.075 1.485 ;
      RECT  14.745 1.485 15.08 1.49 ;
      RECT  14.75 1.49 15.085 1.495 ;
      RECT  14.755 1.495 15.09 1.5 ;
      RECT  14.76 1.5 15.095 1.505 ;
      RECT  14.765 1.505 15.1 1.51 ;
      RECT  14.77 1.51 15.105 1.515 ;
      RECT  14.775 1.515 15.11 1.52 ;
      RECT  14.78 1.52 15.115 1.525 ;
      RECT  14.785 1.525 15.12 1.53 ;
      RECT  14.79 1.53 15.125 1.535 ;
      RECT  14.795 1.535 15.13 1.54 ;
      RECT  14.8 1.54 15.135 1.545 ;
      RECT  14.805 1.545 15.14 1.55 ;
      RECT  14.81 1.55 15.145 1.555 ;
      RECT  14.815 1.555 15.15 1.56 ;
      RECT  14.82 1.56 15.155 1.565 ;
      RECT  14.825 1.565 16.2 1.57 ;
      RECT  14.83 1.57 16.2 1.575 ;
      RECT  14.835 1.575 16.2 1.58 ;
      RECT  14.84 1.58 16.2 1.585 ;
      RECT  14.845 1.585 16.2 1.59 ;
      RECT  14.85 1.59 16.2 1.595 ;
      RECT  14.855 1.595 16.2 1.6 ;
      RECT  14.86 1.6 16.2 1.605 ;
      RECT  14.865 1.605 16.2 1.61 ;
      RECT  14.87 1.61 16.2 1.615 ;
      RECT  14.875 1.615 16.2 1.62 ;
      RECT  14.88 1.62 16.2 1.625 ;
      RECT  14.885 1.625 16.2 1.63 ;
      RECT  14.89 1.63 16.2 1.635 ;
      RECT  14.895 1.635 16.2 1.64 ;
      RECT  14.9 1.64 16.2 1.645 ;
      RECT  14.905 1.645 16.2 1.65 ;
      RECT  14.91 1.65 16.2 1.655 ;
      RECT  14.915 1.655 16.2 1.66 ;
      RECT  14.92 1.66 16.2 1.665 ;
      RECT  14.925 1.665 16.2 1.67 ;
      RECT  14.93 1.67 16.2 1.675 ;
      RECT  14.935 1.675 16.2 1.68 ;
      RECT  14.94 1.68 16.2 1.685 ;
      RECT  14.945 1.685 16.2 1.69 ;
      RECT  14.95 1.69 16.2 1.695 ;
      RECT  14.955 1.695 16.2 1.7 ;
      RECT  14.96 1.7 16.2 1.705 ;
      RECT  14.965 1.705 16.2 1.71 ;
      RECT  14.97 1.71 16.2 1.715 ;
      RECT  14.975 1.715 16.2 1.72 ;
      RECT  14.98 1.72 16.2 1.725 ;
      RECT  14.985 1.725 16.2 1.73 ;
      RECT  14.99 1.73 16.2 1.735 ;
      RECT  14.995 1.735 16.2 1.74 ;
      RECT  15.0 1.74 16.2 1.745 ;
      RECT  15.005 1.745 16.2 1.75 ;
      RECT  15.01 1.75 16.2 1.755 ;
      RECT  15.015 1.755 16.2 1.76 ;
      RECT  15.02 1.76 16.2 1.765 ;
      RECT  15.025 1.765 16.2 1.77 ;
      RECT  15.03 1.77 16.2 1.775 ;
      RECT  15.035 1.775 16.2 1.78 ;
      RECT  15.04 1.78 16.2 1.785 ;
      RECT  15.045 1.785 16.2 1.79 ;
      RECT  15.05 1.79 16.2 1.795 ;
      RECT  3.245 1.005 8.78 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  1.72 1.565 3.475 1.795 ;
      RECT  4.365 1.565 5.0 1.795 ;
      RECT  4.365 1.795 4.595 3.755 ;
      RECT  0.49 3.755 5.0 3.985 ;
      RECT  0.49 3.985 0.72 5.0 ;
      RECT  0.38 5.0 0.72 5.23 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  9.14 1.565 10.195 1.795 ;
      RECT  9.965 1.795 10.195 2.41 ;
      RECT  9.965 2.41 10.68 2.64 ;
      RECT  9.965 2.64 10.195 3.03 ;
      RECT  9.14 3.03 10.195 3.26 ;
      RECT  10.68 1.565 11.315 1.795 ;
      RECT  11.085 1.795 11.315 2.41 ;
      RECT  11.085 2.41 11.93 2.64 ;
      RECT  11.085 2.64 11.315 3.245 ;
      RECT  10.68 3.245 11.315 3.475 ;
      RECT  12.92 1.75 14.675 1.98 ;
      RECT  14.445 1.98 14.675 3.755 ;
      RECT  13.005 3.755 15.5 3.985 ;
      RECT  13.005 3.985 13.235 4.02 ;
      RECT  12.205 4.02 13.235 4.215 ;
      RECT  8.99 4.215 13.235 4.25 ;
      RECT  8.99 4.25 12.435 4.445 ;
      RECT  8.99 4.445 9.22 4.54 ;
      RECT  7.725 4.54 9.22 4.77 ;
      RECT  7.725 4.77 7.955 5.0 ;
      RECT  5.99 5.0 7.955 5.23 ;
      RECT  13.885 2.34 14.115 3.245 ;
      RECT  12.84 3.245 14.115 3.25 ;
      RECT  12.835 3.25 14.115 3.255 ;
      RECT  12.83 3.255 14.115 3.26 ;
      RECT  12.825 3.26 14.115 3.265 ;
      RECT  12.82 3.265 14.115 3.27 ;
      RECT  12.815 3.27 14.115 3.275 ;
      RECT  12.81 3.275 14.115 3.28 ;
      RECT  12.805 3.28 14.115 3.285 ;
      RECT  12.8 3.285 14.115 3.29 ;
      RECT  12.795 3.29 14.115 3.295 ;
      RECT  12.79 3.295 14.115 3.3 ;
      RECT  12.785 3.3 14.115 3.305 ;
      RECT  12.78 3.305 14.115 3.31 ;
      RECT  12.775 3.31 14.115 3.315 ;
      RECT  12.77 3.315 14.115 3.32 ;
      RECT  12.765 3.32 14.115 3.325 ;
      RECT  12.76 3.325 14.115 3.33 ;
      RECT  12.755 3.33 14.115 3.335 ;
      RECT  12.75 3.335 14.115 3.34 ;
      RECT  12.745 3.34 14.115 3.345 ;
      RECT  12.74 3.345 14.115 3.35 ;
      RECT  12.735 3.35 14.115 3.355 ;
      RECT  12.73 3.355 14.115 3.36 ;
      RECT  12.725 3.36 14.115 3.365 ;
      RECT  12.72 3.365 14.115 3.37 ;
      RECT  12.715 3.37 14.115 3.375 ;
      RECT  12.71 3.375 14.115 3.38 ;
      RECT  12.705 3.38 14.115 3.385 ;
      RECT  12.7 3.385 14.115 3.39 ;
      RECT  12.695 3.39 14.115 3.395 ;
      RECT  12.69 3.395 14.115 3.4 ;
      RECT  12.685 3.4 14.115 3.405 ;
      RECT  12.68 3.405 14.115 3.41 ;
      RECT  12.675 3.41 14.115 3.415 ;
      RECT  12.67 3.415 14.115 3.42 ;
      RECT  12.665 3.42 14.115 3.425 ;
      RECT  12.66 3.425 14.115 3.43 ;
      RECT  12.655 3.43 14.115 3.435 ;
      RECT  12.65 3.435 14.115 3.44 ;
      RECT  12.645 3.44 14.115 3.445 ;
      RECT  12.64 3.445 14.115 3.45 ;
      RECT  12.635 3.45 14.115 3.455 ;
      RECT  12.63 3.455 14.115 3.46 ;
      RECT  12.625 3.46 14.115 3.465 ;
      RECT  12.62 3.465 14.115 3.47 ;
      RECT  12.615 3.47 14.115 3.475 ;
      RECT  12.61 3.475 12.935 3.48 ;
      RECT  12.605 3.48 12.93 3.485 ;
      RECT  12.6 3.485 12.925 3.49 ;
      RECT  12.595 3.49 12.92 3.495 ;
      RECT  12.59 3.495 12.915 3.5 ;
      RECT  12.585 3.5 12.91 3.505 ;
      RECT  12.58 3.505 12.905 3.51 ;
      RECT  12.575 3.51 12.9 3.515 ;
      RECT  12.57 3.515 12.895 3.52 ;
      RECT  12.565 3.52 12.89 3.525 ;
      RECT  12.56 3.525 12.885 3.53 ;
      RECT  12.555 3.53 12.88 3.535 ;
      RECT  12.55 3.535 12.875 3.54 ;
      RECT  12.545 3.54 12.87 3.545 ;
      RECT  12.54 3.545 12.865 3.55 ;
      RECT  12.535 3.55 12.86 3.555 ;
      RECT  12.53 3.555 12.855 3.56 ;
      RECT  11.645 3.56 12.85 3.565 ;
      RECT  11.645 3.565 12.845 3.57 ;
      RECT  11.645 3.57 12.84 3.575 ;
      RECT  11.645 3.575 12.835 3.58 ;
      RECT  11.645 3.58 12.83 3.585 ;
      RECT  11.645 3.585 12.825 3.59 ;
      RECT  11.645 3.59 12.82 3.595 ;
      RECT  11.645 3.595 12.815 3.6 ;
      RECT  11.645 3.6 12.81 3.605 ;
      RECT  11.645 3.605 12.805 3.61 ;
      RECT  11.645 3.61 12.8 3.615 ;
      RECT  11.645 3.615 12.795 3.62 ;
      RECT  11.645 3.62 12.79 3.625 ;
      RECT  11.645 3.625 12.785 3.63 ;
      RECT  11.645 3.63 12.78 3.635 ;
      RECT  11.645 3.635 12.775 3.64 ;
      RECT  11.645 3.64 12.77 3.645 ;
      RECT  11.645 3.645 12.765 3.65 ;
      RECT  11.645 3.65 12.76 3.655 ;
      RECT  11.645 3.655 12.755 3.66 ;
      RECT  11.645 3.66 12.75 3.665 ;
      RECT  11.645 3.665 12.745 3.67 ;
      RECT  11.645 3.67 12.74 3.675 ;
      RECT  11.645 3.675 12.735 3.68 ;
      RECT  11.645 3.68 12.73 3.685 ;
      RECT  11.645 3.685 12.725 3.69 ;
      RECT  11.645 3.69 12.72 3.695 ;
      RECT  11.645 3.695 12.715 3.7 ;
      RECT  11.645 3.7 12.71 3.705 ;
      RECT  11.645 3.705 12.705 3.71 ;
      RECT  11.645 3.71 12.7 3.715 ;
      RECT  11.645 3.715 12.695 3.72 ;
      RECT  11.645 3.72 12.69 3.725 ;
      RECT  11.645 3.725 12.685 3.73 ;
      RECT  11.645 3.73 12.68 3.735 ;
      RECT  11.645 3.735 12.675 3.74 ;
      RECT  11.645 3.74 12.67 3.745 ;
      RECT  11.645 3.745 12.665 3.75 ;
      RECT  11.645 3.75 12.66 3.755 ;
      RECT  7.725 1.51 7.955 3.245 ;
      RECT  7.725 3.245 8.8 3.25 ;
      RECT  7.725 3.25 8.805 3.255 ;
      RECT  7.725 3.255 8.81 3.26 ;
      RECT  7.725 3.26 8.815 3.265 ;
      RECT  7.725 3.265 8.82 3.27 ;
      RECT  7.725 3.27 8.825 3.275 ;
      RECT  7.725 3.275 8.83 3.28 ;
      RECT  7.725 3.28 8.835 3.285 ;
      RECT  7.725 3.285 8.84 3.29 ;
      RECT  7.725 3.29 8.845 3.295 ;
      RECT  7.725 3.295 8.85 3.3 ;
      RECT  7.725 3.3 8.855 3.305 ;
      RECT  7.725 3.305 8.86 3.31 ;
      RECT  7.725 3.31 8.865 3.315 ;
      RECT  7.725 3.315 8.87 3.32 ;
      RECT  7.725 3.32 8.875 3.325 ;
      RECT  7.725 3.325 8.88 3.33 ;
      RECT  7.725 3.33 8.885 3.335 ;
      RECT  7.725 3.335 8.89 3.34 ;
      RECT  7.725 3.34 8.895 3.345 ;
      RECT  7.725 3.345 8.9 3.35 ;
      RECT  7.725 3.35 8.905 3.355 ;
      RECT  7.725 3.355 8.91 3.36 ;
      RECT  7.725 3.36 8.915 3.365 ;
      RECT  7.725 3.365 8.92 3.37 ;
      RECT  7.725 3.37 8.925 3.375 ;
      RECT  7.725 3.375 8.93 3.38 ;
      RECT  7.725 3.38 8.935 3.385 ;
      RECT  7.725 3.385 8.94 3.39 ;
      RECT  7.725 3.39 8.945 3.395 ;
      RECT  7.725 3.395 8.95 3.4 ;
      RECT  7.725 3.4 8.955 3.405 ;
      RECT  7.725 3.405 8.96 3.41 ;
      RECT  7.725 3.41 8.965 3.415 ;
      RECT  7.725 3.415 8.97 3.42 ;
      RECT  7.725 3.42 8.975 3.425 ;
      RECT  7.725 3.425 8.98 3.43 ;
      RECT  7.725 3.43 8.985 3.435 ;
      RECT  7.725 3.435 8.99 3.44 ;
      RECT  7.725 3.44 8.995 3.445 ;
      RECT  7.725 3.445 9.0 3.45 ;
      RECT  7.725 3.45 9.005 3.455 ;
      RECT  7.725 3.455 9.01 3.46 ;
      RECT  7.725 3.46 9.015 3.465 ;
      RECT  7.725 3.465 9.02 3.47 ;
      RECT  7.725 3.47 9.025 3.475 ;
      RECT  8.695 3.475 9.03 3.48 ;
      RECT  8.7 3.48 9.035 3.485 ;
      RECT  8.705 3.485 9.04 3.49 ;
      RECT  8.71 3.49 9.045 3.495 ;
      RECT  8.715 3.495 9.05 3.5 ;
      RECT  8.72 3.5 9.055 3.505 ;
      RECT  8.725 3.505 9.06 3.51 ;
      RECT  8.73 3.51 9.065 3.515 ;
      RECT  8.735 3.515 9.07 3.52 ;
      RECT  8.74 3.52 9.075 3.525 ;
      RECT  8.745 3.525 9.08 3.53 ;
      RECT  8.75 3.53 9.085 3.535 ;
      RECT  8.755 3.535 9.09 3.54 ;
      RECT  8.76 3.54 9.095 3.545 ;
      RECT  8.765 3.545 9.1 3.55 ;
      RECT  8.77 3.55 9.105 3.555 ;
      RECT  8.775 3.555 9.11 3.56 ;
      RECT  8.78 3.56 9.115 3.565 ;
      RECT  8.785 3.565 9.12 3.57 ;
      RECT  8.79 3.57 9.125 3.575 ;
      RECT  8.795 3.575 9.13 3.58 ;
      RECT  8.8 3.58 9.135 3.585 ;
      RECT  8.805 3.585 9.14 3.59 ;
      RECT  8.81 3.59 9.145 3.595 ;
      RECT  8.815 3.595 9.15 3.6 ;
      RECT  8.82 3.6 9.155 3.605 ;
      RECT  8.825 3.605 9.16 3.61 ;
      RECT  8.83 3.61 9.165 3.615 ;
      RECT  8.835 3.615 9.17 3.62 ;
      RECT  8.84 3.62 9.175 3.625 ;
      RECT  8.845 3.625 9.18 3.63 ;
      RECT  8.85 3.63 9.185 3.635 ;
      RECT  8.855 3.635 9.19 3.64 ;
      RECT  8.86 3.64 9.195 3.645 ;
      RECT  8.865 3.645 9.2 3.65 ;
      RECT  8.87 3.65 9.205 3.655 ;
      RECT  8.875 3.655 9.21 3.66 ;
      RECT  8.88 3.66 9.215 3.665 ;
      RECT  8.885 3.665 9.22 3.67 ;
      RECT  8.89 3.67 9.225 3.675 ;
      RECT  8.895 3.675 9.23 3.68 ;
      RECT  8.9 3.68 9.235 3.685 ;
      RECT  8.905 3.685 9.24 3.69 ;
      RECT  8.91 3.69 9.245 3.695 ;
      RECT  8.915 3.695 9.25 3.7 ;
      RECT  8.92 3.7 9.255 3.705 ;
      RECT  8.925 3.705 9.26 3.71 ;
      RECT  8.93 3.71 9.265 3.715 ;
      RECT  8.935 3.715 9.27 3.72 ;
      RECT  8.94 3.72 9.275 3.725 ;
      RECT  8.945 3.725 9.28 3.73 ;
      RECT  8.95 3.73 9.285 3.735 ;
      RECT  8.955 3.735 9.29 3.74 ;
      RECT  8.96 3.74 9.295 3.745 ;
      RECT  8.965 3.745 9.3 3.75 ;
      RECT  8.97 3.75 9.305 3.755 ;
      RECT  8.975 3.755 12.655 3.76 ;
      RECT  8.98 3.76 12.65 3.765 ;
      RECT  8.985 3.765 12.645 3.77 ;
      RECT  8.99 3.77 12.64 3.775 ;
      RECT  8.995 3.775 12.635 3.78 ;
      RECT  9.0 3.78 12.63 3.785 ;
      RECT  9.005 3.785 12.625 3.79 ;
      RECT  9.01 3.79 11.875 3.795 ;
      RECT  9.015 3.795 11.875 3.8 ;
      RECT  9.02 3.8 11.875 3.805 ;
      RECT  9.025 3.805 11.875 3.81 ;
      RECT  9.03 3.81 11.875 3.815 ;
      RECT  9.035 3.815 11.875 3.82 ;
      RECT  9.04 3.82 11.875 3.825 ;
      RECT  9.045 3.825 11.875 3.83 ;
      RECT  9.05 3.83 11.875 3.835 ;
      RECT  9.055 3.835 11.875 3.84 ;
      RECT  9.06 3.84 11.875 3.845 ;
      RECT  9.065 3.845 11.875 3.85 ;
      RECT  9.07 3.85 11.875 3.855 ;
      RECT  9.075 3.855 11.875 3.86 ;
      RECT  9.08 3.86 11.875 3.865 ;
      RECT  9.085 3.865 11.875 3.87 ;
      RECT  9.09 3.87 11.875 3.875 ;
      RECT  9.095 3.875 11.875 3.88 ;
      RECT  9.1 3.88 11.875 3.885 ;
      RECT  9.105 3.885 11.875 3.89 ;
      RECT  9.11 3.89 11.875 3.895 ;
      RECT  9.115 3.895 11.875 3.9 ;
      RECT  9.12 3.9 11.875 3.905 ;
      RECT  9.125 3.905 11.875 3.91 ;
      RECT  9.13 3.91 11.875 3.915 ;
      RECT  9.135 3.915 11.875 3.92 ;
      RECT  9.14 3.92 11.875 3.925 ;
      RECT  9.145 3.925 11.875 3.93 ;
      RECT  9.15 3.93 11.875 3.935 ;
      RECT  9.155 3.935 11.875 3.94 ;
      RECT  9.16 3.94 11.875 3.945 ;
      RECT  9.165 3.945 11.875 3.95 ;
      RECT  9.17 3.95 11.875 3.955 ;
      RECT  9.175 3.955 11.875 3.96 ;
      RECT  9.18 3.96 11.875 3.965 ;
      RECT  9.185 3.965 11.875 3.97 ;
      RECT  9.19 3.97 11.875 3.975 ;
      RECT  9.195 3.975 11.875 3.98 ;
      RECT  9.2 3.98 11.875 3.985 ;
      RECT  12.205 1.585 12.435 3.315 ;
      RECT  0.18 3.245 2.76 3.475 ;
      RECT  8.495 3.84 8.725 3.95 ;
      RECT  6.2 3.95 8.725 4.18 ;
      RECT  1.72 4.215 4.3 4.445 ;
      RECT  13.465 4.215 17.74 4.445 ;
      RECT  13.465 4.445 13.695 4.48 ;
      RECT  12.92 4.48 13.695 4.71 ;
      RECT  4.925 4.41 7.24 4.64 ;
      RECT  4.925 4.64 5.155 4.675 ;
      RECT  2.685 4.675 5.155 4.905 ;
      RECT  2.685 4.905 2.915 4.925 ;
      RECT  0.95 4.925 2.915 5.155 ;
      RECT  9.45 4.675 10.71 4.905 ;
      RECT  9.45 4.905 9.68 5.0 ;
      RECT  10.48 4.905 10.71 5.0 ;
      RECT  8.23 5.0 9.68 5.23 ;
      RECT  10.48 5.0 11.92 5.23 ;
      RECT  13.93 4.675 17.48 4.905 ;
      RECT  13.93 4.905 14.16 4.94 ;
      RECT  17.24 4.905 17.48 5.0 ;
      RECT  12.15 4.94 14.16 5.17 ;
      RECT  17.24 5.0 18.65 5.23 ;
  END
END MDN_FSDNSBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDNSBQ_4
#      Description : D-Flip Flop w/scan, neg-edge triggered, lo-async-/set, q-only
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDNSBQ_4
  CLASS CORE ;
  FOREIGN MDN_FSDNSBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 24.64 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 9.635 2.355 ;
      RECT  9.405 2.355 9.635 2.69 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.54 0.6 1.82 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.64 1.565 22.92 1.795 ;
      RECT  22.285 1.795 22.515 3.245 ;
      RECT  19.64 3.245 22.92 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.98 2.12 17.5 2.36 ;
      RECT  14.98 2.36 15.26 2.915 ;
      RECT  17.22 2.36 17.5 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.81 5.74 ;
      RECT  21.165 4.905 21.395 5.46 ;
      RECT  20.72 5.46 21.395 5.74 ;
      RECT  18.925 4.87 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  14.39 5.135 14.73 5.46 ;
      RECT  14.0 5.46 17.36 5.74 ;
      RECT  16.63 5.135 16.97 5.46 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 10.64 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.19 5.135 3.53 5.46 ;
      RECT  2.8 5.46 3.92 5.74 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 24.64 5.74 ;
      LAYER VIA12 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  24.23 5.47 24.49 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 24.81 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  15.12 -0.14 15.85 0.14 ;
      RECT  15.565 0.14 15.795 1.005 ;
      RECT  15.16 1.005 17.74 1.235 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.685 -0.14 3.36 0.14 ;
      RECT  2.685 0.14 2.915 1.005 ;
      RECT  2.42 1.005 2.915 1.23 ;
      RECT  2.42 1.23 2.76 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 24.64 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  22.55 -0.13 22.81 0.13 ;
      RECT  23.11 -0.13 23.37 0.13 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  10.46 0.37 10.81 0.445 ;
      RECT  10.46 0.445 13.05 0.675 ;
      RECT  12.71 0.37 13.05 0.445 ;
      RECT  10.46 0.675 10.69 1.005 ;
      RECT  7.11 0.37 7.45 0.445 ;
      RECT  7.11 0.445 9.635 0.675 ;
      RECT  9.405 0.675 9.635 1.005 ;
      RECT  9.405 1.005 10.69 1.235 ;
      RECT  16.07 0.37 16.41 0.445 ;
      RECT  16.07 0.445 18.33 0.675 ;
      RECT  18.1 0.675 18.33 1.005 ;
      RECT  18.1 1.005 19.155 1.235 ;
      RECT  18.925 1.235 19.155 2.405 ;
      RECT  18.925 2.405 21.825 2.635 ;
      RECT  18.925 2.635 19.155 4.365 ;
      RECT  18.1 4.365 19.155 4.595 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  21.67 0.37 23.13 0.6 ;
      RECT  11.38 1.005 14.605 1.01 ;
      RECT  11.38 1.01 14.61 1.015 ;
      RECT  11.38 1.015 14.615 1.02 ;
      RECT  11.38 1.02 14.62 1.025 ;
      RECT  11.38 1.025 14.625 1.03 ;
      RECT  11.38 1.03 14.63 1.035 ;
      RECT  11.38 1.035 14.635 1.04 ;
      RECT  11.38 1.04 14.64 1.045 ;
      RECT  11.38 1.045 14.645 1.05 ;
      RECT  11.38 1.05 14.65 1.055 ;
      RECT  11.38 1.055 14.655 1.06 ;
      RECT  11.38 1.06 14.66 1.065 ;
      RECT  11.38 1.065 14.665 1.07 ;
      RECT  11.38 1.07 14.67 1.075 ;
      RECT  11.38 1.075 14.675 1.08 ;
      RECT  11.38 1.08 14.68 1.085 ;
      RECT  11.38 1.085 14.685 1.09 ;
      RECT  11.38 1.09 14.69 1.095 ;
      RECT  11.38 1.095 14.695 1.1 ;
      RECT  11.38 1.1 14.7 1.105 ;
      RECT  11.38 1.105 14.705 1.11 ;
      RECT  11.38 1.11 14.71 1.115 ;
      RECT  11.38 1.115 14.715 1.12 ;
      RECT  11.38 1.12 14.72 1.125 ;
      RECT  11.38 1.125 14.725 1.13 ;
      RECT  11.38 1.13 14.73 1.135 ;
      RECT  11.38 1.135 14.735 1.14 ;
      RECT  11.38 1.14 14.74 1.145 ;
      RECT  11.38 1.145 14.745 1.15 ;
      RECT  11.38 1.15 14.75 1.155 ;
      RECT  11.38 1.155 14.755 1.16 ;
      RECT  11.38 1.16 14.76 1.165 ;
      RECT  11.38 1.165 14.765 1.17 ;
      RECT  11.38 1.17 14.77 1.175 ;
      RECT  11.38 1.175 14.775 1.18 ;
      RECT  11.38 1.18 14.78 1.185 ;
      RECT  11.38 1.185 14.785 1.19 ;
      RECT  11.38 1.19 14.79 1.195 ;
      RECT  11.38 1.195 14.795 1.2 ;
      RECT  11.38 1.2 14.8 1.205 ;
      RECT  11.38 1.205 14.805 1.21 ;
      RECT  11.38 1.21 14.81 1.215 ;
      RECT  11.38 1.215 14.815 1.22 ;
      RECT  11.38 1.22 14.82 1.225 ;
      RECT  11.38 1.225 14.825 1.23 ;
      RECT  11.38 1.23 14.83 1.235 ;
      RECT  14.5 1.235 14.835 1.24 ;
      RECT  14.505 1.24 14.84 1.245 ;
      RECT  14.51 1.245 14.845 1.25 ;
      RECT  14.515 1.25 14.85 1.255 ;
      RECT  14.52 1.255 14.855 1.26 ;
      RECT  14.525 1.26 14.86 1.265 ;
      RECT  14.53 1.265 14.865 1.27 ;
      RECT  14.535 1.27 14.87 1.275 ;
      RECT  14.54 1.275 14.875 1.28 ;
      RECT  14.545 1.28 14.88 1.285 ;
      RECT  14.55 1.285 14.885 1.29 ;
      RECT  14.555 1.29 14.89 1.295 ;
      RECT  14.56 1.295 14.895 1.3 ;
      RECT  14.565 1.3 14.9 1.305 ;
      RECT  14.57 1.305 14.905 1.31 ;
      RECT  14.575 1.31 14.91 1.315 ;
      RECT  14.58 1.315 14.915 1.32 ;
      RECT  14.585 1.32 14.92 1.325 ;
      RECT  14.59 1.325 14.925 1.33 ;
      RECT  14.595 1.33 14.93 1.335 ;
      RECT  14.6 1.335 14.935 1.34 ;
      RECT  14.605 1.34 14.94 1.345 ;
      RECT  14.61 1.345 14.945 1.35 ;
      RECT  14.615 1.35 14.95 1.355 ;
      RECT  14.62 1.355 14.955 1.36 ;
      RECT  14.625 1.36 14.96 1.365 ;
      RECT  14.63 1.365 14.965 1.37 ;
      RECT  14.635 1.37 14.97 1.375 ;
      RECT  14.64 1.375 14.975 1.38 ;
      RECT  14.645 1.38 14.98 1.385 ;
      RECT  14.65 1.385 14.985 1.39 ;
      RECT  14.655 1.39 14.99 1.395 ;
      RECT  14.66 1.395 14.995 1.4 ;
      RECT  14.665 1.4 15.0 1.405 ;
      RECT  14.67 1.405 15.005 1.41 ;
      RECT  14.675 1.41 15.01 1.415 ;
      RECT  14.68 1.415 15.015 1.42 ;
      RECT  14.685 1.42 15.02 1.425 ;
      RECT  14.69 1.425 15.025 1.43 ;
      RECT  14.695 1.43 15.03 1.435 ;
      RECT  14.7 1.435 15.035 1.44 ;
      RECT  14.705 1.44 15.04 1.445 ;
      RECT  14.71 1.445 15.045 1.45 ;
      RECT  14.715 1.45 15.05 1.455 ;
      RECT  14.72 1.455 15.055 1.46 ;
      RECT  14.725 1.46 15.06 1.465 ;
      RECT  14.73 1.465 15.065 1.47 ;
      RECT  14.735 1.47 15.07 1.475 ;
      RECT  14.74 1.475 15.075 1.48 ;
      RECT  14.745 1.48 15.08 1.485 ;
      RECT  14.75 1.485 15.085 1.49 ;
      RECT  14.755 1.49 15.09 1.495 ;
      RECT  14.76 1.495 15.095 1.5 ;
      RECT  14.765 1.5 15.1 1.505 ;
      RECT  14.77 1.505 15.105 1.51 ;
      RECT  14.775 1.51 15.11 1.515 ;
      RECT  14.78 1.515 15.115 1.52 ;
      RECT  14.785 1.52 15.12 1.525 ;
      RECT  14.79 1.525 15.125 1.53 ;
      RECT  14.795 1.53 15.13 1.535 ;
      RECT  14.8 1.535 15.135 1.54 ;
      RECT  14.805 1.54 15.14 1.545 ;
      RECT  14.81 1.545 15.145 1.55 ;
      RECT  14.815 1.55 15.15 1.555 ;
      RECT  14.82 1.555 15.155 1.56 ;
      RECT  14.825 1.56 15.16 1.565 ;
      RECT  14.83 1.565 16.205 1.57 ;
      RECT  14.835 1.57 16.205 1.575 ;
      RECT  14.84 1.575 16.205 1.58 ;
      RECT  14.845 1.58 16.205 1.585 ;
      RECT  14.85 1.585 16.205 1.59 ;
      RECT  14.855 1.59 16.205 1.595 ;
      RECT  14.86 1.595 16.205 1.6 ;
      RECT  14.865 1.6 16.205 1.605 ;
      RECT  14.87 1.605 16.205 1.61 ;
      RECT  14.875 1.61 16.205 1.615 ;
      RECT  14.88 1.615 16.205 1.62 ;
      RECT  14.885 1.62 16.205 1.625 ;
      RECT  14.89 1.625 16.205 1.63 ;
      RECT  14.895 1.63 16.205 1.635 ;
      RECT  14.9 1.635 16.205 1.64 ;
      RECT  14.905 1.64 16.205 1.645 ;
      RECT  14.91 1.645 16.205 1.65 ;
      RECT  14.915 1.65 16.205 1.655 ;
      RECT  14.92 1.655 16.205 1.66 ;
      RECT  14.925 1.66 16.205 1.665 ;
      RECT  14.93 1.665 16.205 1.67 ;
      RECT  14.935 1.67 16.205 1.675 ;
      RECT  14.94 1.675 16.205 1.68 ;
      RECT  14.945 1.68 16.205 1.685 ;
      RECT  14.95 1.685 16.205 1.69 ;
      RECT  14.955 1.69 16.205 1.695 ;
      RECT  14.96 1.695 16.205 1.7 ;
      RECT  14.965 1.7 16.205 1.705 ;
      RECT  14.97 1.705 16.205 1.71 ;
      RECT  14.975 1.71 16.205 1.715 ;
      RECT  14.98 1.715 16.205 1.72 ;
      RECT  14.985 1.72 16.205 1.725 ;
      RECT  14.99 1.725 16.205 1.73 ;
      RECT  14.995 1.73 16.205 1.735 ;
      RECT  15.0 1.735 16.205 1.74 ;
      RECT  15.005 1.74 16.205 1.745 ;
      RECT  15.01 1.745 16.205 1.75 ;
      RECT  15.015 1.75 16.205 1.755 ;
      RECT  15.02 1.755 16.205 1.76 ;
      RECT  15.025 1.76 16.205 1.765 ;
      RECT  15.03 1.765 16.205 1.77 ;
      RECT  15.035 1.77 16.205 1.775 ;
      RECT  15.04 1.775 16.205 1.78 ;
      RECT  15.045 1.78 16.205 1.785 ;
      RECT  15.05 1.785 16.205 1.79 ;
      RECT  15.055 1.79 16.205 1.795 ;
      RECT  3.245 1.005 8.78 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  1.72 1.565 3.475 1.795 ;
      RECT  12.92 1.565 14.27 1.57 ;
      RECT  12.92 1.57 14.275 1.575 ;
      RECT  12.92 1.575 14.28 1.58 ;
      RECT  12.92 1.58 14.285 1.585 ;
      RECT  12.92 1.585 14.29 1.59 ;
      RECT  12.92 1.59 14.295 1.595 ;
      RECT  12.92 1.595 14.3 1.6 ;
      RECT  12.92 1.6 14.305 1.605 ;
      RECT  12.92 1.605 14.31 1.61 ;
      RECT  12.92 1.61 14.315 1.615 ;
      RECT  12.92 1.615 14.32 1.62 ;
      RECT  12.92 1.62 14.325 1.625 ;
      RECT  12.92 1.625 14.33 1.63 ;
      RECT  12.92 1.63 14.335 1.635 ;
      RECT  12.92 1.635 14.34 1.64 ;
      RECT  12.92 1.64 14.345 1.645 ;
      RECT  12.92 1.645 14.35 1.65 ;
      RECT  12.92 1.65 14.355 1.655 ;
      RECT  12.92 1.655 14.36 1.66 ;
      RECT  12.92 1.66 14.365 1.665 ;
      RECT  12.92 1.665 14.37 1.67 ;
      RECT  12.92 1.67 14.375 1.675 ;
      RECT  12.92 1.675 14.38 1.68 ;
      RECT  12.92 1.68 14.385 1.685 ;
      RECT  12.92 1.685 14.39 1.69 ;
      RECT  12.92 1.69 14.395 1.695 ;
      RECT  12.92 1.695 14.4 1.7 ;
      RECT  12.92 1.7 14.405 1.705 ;
      RECT  12.92 1.705 14.41 1.71 ;
      RECT  12.92 1.71 14.415 1.715 ;
      RECT  12.92 1.715 14.42 1.72 ;
      RECT  12.92 1.72 14.425 1.725 ;
      RECT  12.92 1.725 14.43 1.73 ;
      RECT  12.92 1.73 14.435 1.735 ;
      RECT  12.92 1.735 14.44 1.74 ;
      RECT  12.92 1.74 14.445 1.745 ;
      RECT  12.92 1.745 14.45 1.75 ;
      RECT  12.92 1.75 14.455 1.755 ;
      RECT  12.92 1.755 14.46 1.76 ;
      RECT  12.92 1.76 14.465 1.765 ;
      RECT  12.92 1.765 14.47 1.77 ;
      RECT  12.92 1.77 14.475 1.775 ;
      RECT  12.92 1.775 14.48 1.78 ;
      RECT  12.92 1.78 14.485 1.785 ;
      RECT  12.92 1.785 14.49 1.79 ;
      RECT  12.92 1.79 14.495 1.795 ;
      RECT  14.165 1.795 14.5 1.8 ;
      RECT  14.17 1.8 14.505 1.805 ;
      RECT  14.175 1.805 14.51 1.81 ;
      RECT  14.18 1.81 14.515 1.815 ;
      RECT  14.185 1.815 14.52 1.82 ;
      RECT  14.19 1.82 14.525 1.825 ;
      RECT  14.195 1.825 14.53 1.83 ;
      RECT  14.2 1.83 14.535 1.835 ;
      RECT  14.205 1.835 14.54 1.84 ;
      RECT  14.21 1.84 14.545 1.845 ;
      RECT  14.215 1.845 14.55 1.85 ;
      RECT  14.22 1.85 14.555 1.855 ;
      RECT  14.225 1.855 14.56 1.86 ;
      RECT  14.23 1.86 14.565 1.865 ;
      RECT  14.235 1.865 14.57 1.87 ;
      RECT  14.24 1.87 14.575 1.875 ;
      RECT  14.245 1.875 14.58 1.88 ;
      RECT  14.25 1.88 14.585 1.885 ;
      RECT  14.255 1.885 14.59 1.89 ;
      RECT  14.26 1.89 14.595 1.895 ;
      RECT  14.265 1.895 14.6 1.9 ;
      RECT  14.27 1.9 14.605 1.905 ;
      RECT  14.275 1.905 14.61 1.91 ;
      RECT  14.28 1.91 14.615 1.915 ;
      RECT  14.285 1.915 14.62 1.92 ;
      RECT  14.29 1.92 14.625 1.925 ;
      RECT  14.295 1.925 14.63 1.93 ;
      RECT  14.3 1.93 14.635 1.935 ;
      RECT  14.305 1.935 14.64 1.94 ;
      RECT  14.31 1.94 14.645 1.945 ;
      RECT  14.315 1.945 14.65 1.95 ;
      RECT  14.32 1.95 14.655 1.955 ;
      RECT  14.325 1.955 14.66 1.96 ;
      RECT  14.33 1.96 14.665 1.965 ;
      RECT  14.335 1.965 14.67 1.97 ;
      RECT  14.34 1.97 14.675 1.975 ;
      RECT  14.345 1.975 14.675 1.98 ;
      RECT  14.35 1.98 14.675 1.985 ;
      RECT  14.355 1.985 14.675 1.99 ;
      RECT  14.36 1.99 14.675 1.995 ;
      RECT  14.365 1.995 14.675 2.0 ;
      RECT  14.37 2.0 14.675 2.005 ;
      RECT  14.375 2.005 14.675 2.01 ;
      RECT  14.38 2.01 14.675 2.015 ;
      RECT  14.385 2.015 14.675 2.02 ;
      RECT  14.39 2.02 14.675 2.025 ;
      RECT  14.395 2.025 14.675 2.03 ;
      RECT  14.4 2.03 14.675 2.035 ;
      RECT  14.405 2.035 14.675 2.04 ;
      RECT  14.41 2.04 14.675 2.045 ;
      RECT  14.415 2.045 14.675 2.05 ;
      RECT  14.42 2.05 14.675 2.055 ;
      RECT  14.425 2.055 14.675 2.06 ;
      RECT  14.43 2.06 14.675 2.065 ;
      RECT  14.435 2.065 14.675 2.07 ;
      RECT  14.44 2.07 14.675 2.075 ;
      RECT  14.445 2.075 14.675 3.75 ;
      RECT  13.01 3.75 15.5 3.98 ;
      RECT  13.01 3.98 13.24 4.01 ;
      RECT  12.205 4.01 13.24 4.24 ;
      RECT  12.205 4.24 12.435 4.365 ;
      RECT  8.98 4.205 11.315 4.365 ;
      RECT  8.98 4.365 12.435 4.435 ;
      RECT  8.98 4.435 9.21 4.54 ;
      RECT  11.085 4.435 12.435 4.595 ;
      RECT  7.725 4.54 9.21 4.77 ;
      RECT  7.725 4.77 7.955 5.0 ;
      RECT  5.99 5.0 7.955 5.23 ;
      RECT  4.365 1.565 5.0 1.795 ;
      RECT  4.365 1.795 4.595 3.755 ;
      RECT  0.49 3.755 5.0 3.985 ;
      RECT  0.49 3.985 0.72 5.0 ;
      RECT  0.38 5.0 0.72 5.23 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  9.14 1.565 10.195 1.795 ;
      RECT  9.965 1.795 10.195 2.405 ;
      RECT  9.965 2.405 10.81 2.635 ;
      RECT  9.965 2.635 10.195 3.03 ;
      RECT  9.14 3.03 10.195 3.26 ;
      RECT  10.68 1.565 11.315 1.795 ;
      RECT  11.085 1.795 11.315 2.405 ;
      RECT  11.085 2.405 11.93 2.635 ;
      RECT  11.085 2.635 11.315 3.245 ;
      RECT  10.68 3.245 11.315 3.475 ;
      RECT  13.885 2.365 14.115 3.245 ;
      RECT  12.85 3.245 14.115 3.25 ;
      RECT  12.845 3.25 14.115 3.255 ;
      RECT  12.84 3.255 14.115 3.26 ;
      RECT  12.835 3.26 14.115 3.265 ;
      RECT  12.83 3.265 14.115 3.27 ;
      RECT  12.825 3.27 14.115 3.275 ;
      RECT  12.82 3.275 14.115 3.28 ;
      RECT  12.815 3.28 14.115 3.285 ;
      RECT  12.81 3.285 14.115 3.29 ;
      RECT  12.805 3.29 14.115 3.295 ;
      RECT  12.8 3.295 14.115 3.3 ;
      RECT  12.795 3.3 14.115 3.305 ;
      RECT  12.79 3.305 14.115 3.31 ;
      RECT  12.785 3.31 14.115 3.315 ;
      RECT  12.78 3.315 14.115 3.32 ;
      RECT  12.775 3.32 14.115 3.325 ;
      RECT  12.77 3.325 14.115 3.33 ;
      RECT  12.765 3.33 14.115 3.335 ;
      RECT  12.76 3.335 14.115 3.34 ;
      RECT  12.755 3.34 14.115 3.345 ;
      RECT  12.75 3.345 14.115 3.35 ;
      RECT  12.745 3.35 14.115 3.355 ;
      RECT  12.74 3.355 14.115 3.36 ;
      RECT  12.735 3.36 14.115 3.365 ;
      RECT  12.73 3.365 14.115 3.37 ;
      RECT  12.725 3.37 14.115 3.375 ;
      RECT  12.72 3.375 14.115 3.38 ;
      RECT  12.715 3.38 14.115 3.385 ;
      RECT  12.71 3.385 14.115 3.39 ;
      RECT  12.705 3.39 14.115 3.395 ;
      RECT  12.7 3.395 14.115 3.4 ;
      RECT  12.695 3.4 14.115 3.405 ;
      RECT  12.69 3.405 14.115 3.41 ;
      RECT  12.685 3.41 14.115 3.415 ;
      RECT  12.68 3.415 14.115 3.42 ;
      RECT  12.675 3.42 14.115 3.425 ;
      RECT  12.67 3.425 14.115 3.43 ;
      RECT  12.665 3.43 14.115 3.435 ;
      RECT  12.66 3.435 14.115 3.44 ;
      RECT  12.655 3.44 14.115 3.445 ;
      RECT  12.65 3.445 14.115 3.45 ;
      RECT  12.645 3.45 14.115 3.455 ;
      RECT  12.64 3.455 14.115 3.46 ;
      RECT  12.635 3.46 14.115 3.465 ;
      RECT  12.63 3.465 14.115 3.47 ;
      RECT  12.625 3.47 14.11 3.475 ;
      RECT  12.62 3.475 12.945 3.48 ;
      RECT  12.615 3.48 12.94 3.485 ;
      RECT  12.61 3.485 12.935 3.49 ;
      RECT  12.605 3.49 12.93 3.495 ;
      RECT  12.6 3.495 12.925 3.5 ;
      RECT  12.595 3.5 12.92 3.505 ;
      RECT  12.59 3.505 12.915 3.51 ;
      RECT  12.585 3.51 12.91 3.515 ;
      RECT  12.58 3.515 12.905 3.52 ;
      RECT  12.575 3.52 12.9 3.525 ;
      RECT  12.57 3.525 12.895 3.53 ;
      RECT  12.565 3.53 12.89 3.535 ;
      RECT  12.56 3.535 12.885 3.54 ;
      RECT  12.555 3.54 12.88 3.545 ;
      RECT  12.55 3.545 12.875 3.55 ;
      RECT  11.645 3.55 12.87 3.555 ;
      RECT  11.645 3.555 12.865 3.56 ;
      RECT  11.645 3.56 12.86 3.565 ;
      RECT  11.645 3.565 12.855 3.57 ;
      RECT  11.645 3.57 12.85 3.575 ;
      RECT  11.645 3.575 12.845 3.58 ;
      RECT  11.645 3.58 12.84 3.585 ;
      RECT  11.645 3.585 12.835 3.59 ;
      RECT  11.645 3.59 12.83 3.595 ;
      RECT  11.645 3.595 12.825 3.6 ;
      RECT  11.645 3.6 12.82 3.605 ;
      RECT  11.645 3.605 12.815 3.61 ;
      RECT  11.645 3.61 12.81 3.615 ;
      RECT  11.645 3.615 12.805 3.62 ;
      RECT  11.645 3.62 12.8 3.625 ;
      RECT  11.645 3.625 12.795 3.63 ;
      RECT  11.645 3.63 12.79 3.635 ;
      RECT  11.645 3.635 12.785 3.64 ;
      RECT  11.645 3.64 12.78 3.645 ;
      RECT  11.645 3.645 12.775 3.65 ;
      RECT  11.645 3.65 12.77 3.655 ;
      RECT  11.645 3.655 12.765 3.66 ;
      RECT  11.645 3.66 12.76 3.665 ;
      RECT  11.645 3.665 12.755 3.67 ;
      RECT  11.645 3.67 12.75 3.675 ;
      RECT  11.645 3.675 12.745 3.68 ;
      RECT  11.645 3.68 12.74 3.685 ;
      RECT  11.645 3.685 12.735 3.69 ;
      RECT  11.645 3.69 12.73 3.695 ;
      RECT  11.645 3.695 12.725 3.7 ;
      RECT  11.645 3.7 12.72 3.705 ;
      RECT  11.645 3.705 12.715 3.71 ;
      RECT  11.645 3.71 12.71 3.715 ;
      RECT  11.645 3.715 12.705 3.72 ;
      RECT  11.645 3.72 12.7 3.725 ;
      RECT  11.645 3.725 12.695 3.73 ;
      RECT  11.645 3.73 12.69 3.735 ;
      RECT  11.645 3.735 12.685 3.74 ;
      RECT  11.645 3.74 12.68 3.745 ;
      RECT  7.725 1.51 7.955 3.245 ;
      RECT  7.725 3.245 8.74 3.25 ;
      RECT  7.725 3.25 8.745 3.255 ;
      RECT  7.725 3.255 8.75 3.26 ;
      RECT  7.725 3.26 8.755 3.265 ;
      RECT  7.725 3.265 8.76 3.27 ;
      RECT  7.725 3.27 8.765 3.275 ;
      RECT  7.725 3.275 8.77 3.28 ;
      RECT  7.725 3.28 8.775 3.285 ;
      RECT  7.725 3.285 8.78 3.29 ;
      RECT  7.725 3.29 8.785 3.295 ;
      RECT  7.725 3.295 8.79 3.3 ;
      RECT  7.725 3.3 8.795 3.305 ;
      RECT  7.725 3.305 8.8 3.31 ;
      RECT  7.725 3.31 8.805 3.315 ;
      RECT  7.725 3.315 8.81 3.32 ;
      RECT  7.725 3.32 8.815 3.325 ;
      RECT  7.725 3.325 8.82 3.33 ;
      RECT  7.725 3.33 8.825 3.335 ;
      RECT  7.725 3.335 8.83 3.34 ;
      RECT  7.725 3.34 8.835 3.345 ;
      RECT  7.725 3.345 8.84 3.35 ;
      RECT  7.725 3.35 8.845 3.355 ;
      RECT  7.725 3.355 8.85 3.36 ;
      RECT  7.725 3.36 8.855 3.365 ;
      RECT  7.725 3.365 8.86 3.37 ;
      RECT  7.725 3.37 8.865 3.375 ;
      RECT  7.725 3.375 8.87 3.38 ;
      RECT  7.725 3.38 8.875 3.385 ;
      RECT  7.725 3.385 8.88 3.39 ;
      RECT  7.725 3.39 8.885 3.395 ;
      RECT  7.725 3.395 8.89 3.4 ;
      RECT  7.725 3.4 8.895 3.405 ;
      RECT  7.725 3.405 8.9 3.41 ;
      RECT  7.725 3.41 8.905 3.415 ;
      RECT  7.725 3.415 8.91 3.42 ;
      RECT  7.725 3.42 8.915 3.425 ;
      RECT  7.725 3.425 8.92 3.43 ;
      RECT  7.725 3.43 8.925 3.435 ;
      RECT  7.725 3.435 8.93 3.44 ;
      RECT  7.725 3.44 8.935 3.445 ;
      RECT  7.725 3.445 8.94 3.45 ;
      RECT  7.725 3.45 8.945 3.455 ;
      RECT  7.725 3.455 8.95 3.46 ;
      RECT  7.725 3.46 8.955 3.465 ;
      RECT  7.725 3.465 8.96 3.47 ;
      RECT  7.725 3.47 8.965 3.475 ;
      RECT  8.635 3.475 8.97 3.48 ;
      RECT  8.64 3.48 8.975 3.485 ;
      RECT  8.645 3.485 8.98 3.49 ;
      RECT  8.65 3.49 8.985 3.495 ;
      RECT  8.655 3.495 8.99 3.5 ;
      RECT  8.66 3.5 8.995 3.505 ;
      RECT  8.665 3.505 9.0 3.51 ;
      RECT  8.67 3.51 9.005 3.515 ;
      RECT  8.675 3.515 9.01 3.52 ;
      RECT  8.68 3.52 9.015 3.525 ;
      RECT  8.685 3.525 9.02 3.53 ;
      RECT  8.69 3.53 9.025 3.535 ;
      RECT  8.695 3.535 9.03 3.54 ;
      RECT  8.7 3.54 9.035 3.545 ;
      RECT  8.705 3.545 9.04 3.55 ;
      RECT  8.71 3.55 9.045 3.555 ;
      RECT  8.715 3.555 9.05 3.56 ;
      RECT  8.72 3.56 9.055 3.565 ;
      RECT  8.725 3.565 9.06 3.57 ;
      RECT  8.73 3.57 9.065 3.575 ;
      RECT  8.735 3.575 9.07 3.58 ;
      RECT  8.74 3.58 9.075 3.585 ;
      RECT  8.745 3.585 9.08 3.59 ;
      RECT  8.75 3.59 9.085 3.595 ;
      RECT  8.755 3.595 9.09 3.6 ;
      RECT  8.76 3.6 9.095 3.605 ;
      RECT  8.765 3.605 9.1 3.61 ;
      RECT  8.77 3.61 9.105 3.615 ;
      RECT  8.775 3.615 9.11 3.62 ;
      RECT  8.78 3.62 9.115 3.625 ;
      RECT  8.785 3.625 9.12 3.63 ;
      RECT  8.79 3.63 9.125 3.635 ;
      RECT  8.795 3.635 9.13 3.64 ;
      RECT  8.8 3.64 9.135 3.645 ;
      RECT  8.805 3.645 9.14 3.65 ;
      RECT  8.81 3.65 9.145 3.655 ;
      RECT  8.815 3.655 9.15 3.66 ;
      RECT  8.82 3.66 9.155 3.665 ;
      RECT  8.825 3.665 9.16 3.67 ;
      RECT  8.83 3.67 9.165 3.675 ;
      RECT  8.835 3.675 9.17 3.68 ;
      RECT  8.84 3.68 9.175 3.685 ;
      RECT  8.845 3.685 9.18 3.69 ;
      RECT  8.85 3.69 9.185 3.695 ;
      RECT  8.855 3.695 9.19 3.7 ;
      RECT  8.86 3.7 9.195 3.705 ;
      RECT  8.865 3.705 9.2 3.71 ;
      RECT  8.87 3.71 9.205 3.715 ;
      RECT  8.875 3.715 9.21 3.72 ;
      RECT  8.88 3.72 9.215 3.725 ;
      RECT  8.885 3.725 9.22 3.73 ;
      RECT  8.89 3.73 9.225 3.735 ;
      RECT  8.895 3.735 9.23 3.74 ;
      RECT  8.9 3.74 9.235 3.745 ;
      RECT  8.905 3.745 12.675 3.75 ;
      RECT  8.91 3.75 12.67 3.755 ;
      RECT  8.915 3.755 12.665 3.76 ;
      RECT  8.92 3.76 12.66 3.765 ;
      RECT  8.925 3.765 12.655 3.77 ;
      RECT  8.93 3.77 12.65 3.775 ;
      RECT  8.935 3.775 12.645 3.78 ;
      RECT  8.94 3.78 11.875 3.785 ;
      RECT  8.945 3.785 11.875 3.79 ;
      RECT  8.95 3.79 11.875 3.795 ;
      RECT  8.955 3.795 11.875 3.8 ;
      RECT  8.96 3.8 11.875 3.805 ;
      RECT  8.965 3.805 11.875 3.81 ;
      RECT  8.97 3.81 11.875 3.815 ;
      RECT  8.975 3.815 11.875 3.82 ;
      RECT  8.98 3.82 11.875 3.825 ;
      RECT  8.985 3.825 11.875 3.83 ;
      RECT  8.99 3.83 11.875 3.835 ;
      RECT  8.995 3.835 11.875 3.84 ;
      RECT  9.0 3.84 11.875 3.845 ;
      RECT  9.005 3.845 11.875 3.85 ;
      RECT  9.01 3.85 11.875 3.855 ;
      RECT  9.015 3.855 11.875 3.86 ;
      RECT  9.02 3.86 11.875 3.865 ;
      RECT  9.025 3.865 11.875 3.87 ;
      RECT  9.03 3.87 11.875 3.875 ;
      RECT  9.035 3.875 11.875 3.88 ;
      RECT  9.04 3.88 11.875 3.885 ;
      RECT  9.045 3.885 11.875 3.89 ;
      RECT  9.05 3.89 11.875 3.895 ;
      RECT  9.055 3.895 11.875 3.9 ;
      RECT  9.06 3.9 11.875 3.905 ;
      RECT  9.065 3.905 11.875 3.91 ;
      RECT  9.07 3.91 11.875 3.915 ;
      RECT  9.075 3.915 11.875 3.92 ;
      RECT  9.08 3.92 11.875 3.925 ;
      RECT  9.085 3.925 11.875 3.93 ;
      RECT  9.09 3.93 11.875 3.935 ;
      RECT  9.095 3.935 11.875 3.94 ;
      RECT  9.1 3.94 11.875 3.945 ;
      RECT  9.105 3.945 11.875 3.95 ;
      RECT  9.11 3.95 11.875 3.955 ;
      RECT  9.115 3.955 11.875 3.96 ;
      RECT  9.12 3.96 11.875 3.965 ;
      RECT  9.125 3.965 11.875 3.97 ;
      RECT  9.13 3.97 11.875 3.975 ;
      RECT  12.205 1.51 12.435 3.315 ;
      RECT  0.18 3.245 2.76 3.475 ;
      RECT  6.2 3.935 8.725 4.165 ;
      RECT  8.495 4.165 8.725 4.275 ;
      RECT  1.72 4.215 4.3 4.445 ;
      RECT  13.47 4.215 17.74 4.445 ;
      RECT  13.47 4.445 13.7 4.48 ;
      RECT  12.92 4.48 13.7 4.71 ;
      RECT  4.925 4.41 7.24 4.64 ;
      RECT  4.925 4.64 5.155 4.675 ;
      RECT  2.685 4.675 5.155 4.905 ;
      RECT  2.685 4.905 2.915 4.925 ;
      RECT  0.95 4.925 2.915 5.155 ;
      RECT  9.44 4.665 10.755 4.905 ;
      RECT  9.44 4.905 9.68 5.0 ;
      RECT  10.525 4.905 10.755 5.0 ;
      RECT  8.23 5.0 9.68 5.23 ;
      RECT  10.525 5.0 11.92 5.23 ;
      RECT  13.93 4.675 17.475 4.905 ;
      RECT  13.93 4.905 14.16 4.985 ;
      RECT  17.245 4.905 17.475 5.0 ;
      RECT  12.15 4.985 14.16 5.215 ;
      RECT  17.245 5.0 18.65 5.23 ;
  END
END MDN_FSDNSBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDP_4
#      Description : D-Flip Flop w/scan, pos-edge triggered
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDP_4
  CLASS CORE ;
  FOREIGN MDN_FSDP_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 26.88 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.4 1.565 21.395 1.795 ;
      RECT  21.165 1.795 21.395 3.245 ;
      RECT  17.4 3.245 21.395 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  22.58 1.565 26.7 1.795 ;
      RECT  24.525 1.795 24.755 3.245 ;
      RECT  22.58 3.245 26.7 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.645 5.46 27.05 5.74 ;
      RECT  23.405 4.905 23.635 5.46 ;
      RECT  23.405 5.46 24.08 5.74 ;
      RECT  21.165 4.905 21.395 5.46 ;
      RECT  21.165 5.46 21.84 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 12.435 5.74 ;
      RECT  12.205 5.0 12.435 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 26.88 5.74 ;
      LAYER VIA12 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 -0.14 27.05 0.14 ;
      RECT  25.645 0.14 25.875 0.7 ;
      RECT  23.405 -0.14 24.08 0.14 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  21.165 -0.14 21.84 0.14 ;
      RECT  21.165 0.14 21.395 0.73 ;
      RECT  18.925 -0.14 19.6 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  3.805 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.805 0.14 4.035 0.89 ;
      RECT  3.805 0.89 4.3 1.12 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 26.88 0.14 ;
      LAYER VIA12 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.46 0.6 ;
      RECT  6.23 0.6 6.46 0.83 ;
      RECT  6.23 0.83 9.635 1.005 ;
      RECT  6.23 1.005 12.435 1.06 ;
      RECT  9.41 1.06 12.435 1.235 ;
      RECT  12.205 1.235 12.435 1.75 ;
      RECT  12.205 1.75 13.96 1.98 ;
      RECT  12.205 1.98 12.435 3.245 ;
      RECT  11.38 3.245 12.435 3.475 ;
      RECT  12.205 3.475 12.435 3.62 ;
      RECT  12.205 3.62 14.115 3.805 ;
      RECT  12.205 3.805 15.5 3.85 ;
      RECT  13.885 3.85 15.5 4.035 ;
      RECT  7.11 0.37 9.69 0.6 ;
      RECT  12.71 0.37 13.225 0.6 ;
      RECT  12.995 0.6 13.225 0.83 ;
      RECT  12.995 0.83 16.09 1.06 ;
      RECT  15.86 1.06 16.09 1.565 ;
      RECT  15.86 1.565 16.355 1.795 ;
      RECT  16.125 1.795 16.355 2.125 ;
      RECT  16.125 2.125 20.835 2.355 ;
      RECT  17.245 2.355 17.475 2.69 ;
      RECT  18.365 2.355 18.595 2.69 ;
      RECT  19.485 2.355 19.715 2.69 ;
      RECT  20.605 2.355 20.835 2.69 ;
      RECT  16.125 2.355 16.355 3.245 ;
      RECT  15.86 3.245 16.355 3.475 ;
      RECT  14.39 0.37 16.41 0.6 ;
      RECT  21.67 0.37 22.01 0.6 ;
      RECT  21.67 0.6 21.9 1.005 ;
      RECT  20.55 0.37 20.89 0.6 ;
      RECT  20.66 0.6 20.89 1.005 ;
      RECT  20.66 1.005 21.9 1.235 ;
      RECT  23.91 0.37 25.37 0.6 ;
      RECT  4.75 1.005 5.715 1.01 ;
      RECT  4.745 1.01 5.715 1.015 ;
      RECT  4.74 1.015 5.715 1.02 ;
      RECT  4.735 1.02 5.715 1.025 ;
      RECT  4.73 1.025 5.715 1.03 ;
      RECT  4.725 1.03 5.715 1.035 ;
      RECT  4.72 1.035 5.715 1.04 ;
      RECT  4.715 1.04 5.715 1.045 ;
      RECT  4.71 1.045 5.715 1.05 ;
      RECT  4.705 1.05 5.715 1.055 ;
      RECT  4.7 1.055 5.715 1.06 ;
      RECT  4.695 1.06 5.715 1.065 ;
      RECT  4.69 1.065 5.715 1.07 ;
      RECT  4.685 1.07 5.715 1.075 ;
      RECT  4.68 1.075 5.715 1.08 ;
      RECT  4.675 1.08 5.715 1.085 ;
      RECT  4.67 1.085 5.715 1.09 ;
      RECT  4.665 1.09 5.715 1.095 ;
      RECT  4.66 1.095 5.715 1.1 ;
      RECT  4.655 1.1 5.715 1.105 ;
      RECT  4.65 1.105 5.715 1.11 ;
      RECT  4.645 1.11 5.715 1.115 ;
      RECT  4.64 1.115 5.715 1.12 ;
      RECT  4.635 1.12 5.715 1.125 ;
      RECT  4.63 1.125 5.715 1.13 ;
      RECT  4.625 1.13 5.715 1.135 ;
      RECT  4.62 1.135 5.715 1.14 ;
      RECT  4.615 1.14 5.715 1.145 ;
      RECT  4.61 1.145 5.715 1.15 ;
      RECT  4.605 1.15 5.715 1.155 ;
      RECT  4.6 1.155 5.715 1.16 ;
      RECT  4.595 1.16 5.715 1.165 ;
      RECT  4.59 1.165 5.715 1.17 ;
      RECT  4.585 1.17 5.715 1.175 ;
      RECT  4.58 1.175 5.715 1.18 ;
      RECT  4.575 1.18 5.715 1.185 ;
      RECT  4.57 1.185 5.715 1.19 ;
      RECT  4.565 1.19 5.715 1.195 ;
      RECT  4.56 1.195 5.715 1.2 ;
      RECT  4.555 1.2 5.715 1.205 ;
      RECT  4.55 1.205 5.715 1.21 ;
      RECT  4.545 1.21 5.715 1.215 ;
      RECT  4.54 1.215 5.715 1.22 ;
      RECT  4.535 1.22 5.715 1.225 ;
      RECT  4.53 1.225 5.715 1.23 ;
      RECT  4.525 1.23 5.715 1.235 ;
      RECT  4.52 1.235 4.845 1.24 ;
      RECT  5.485 1.235 5.715 1.75 ;
      RECT  4.515 1.24 4.84 1.245 ;
      RECT  4.51 1.245 4.835 1.25 ;
      RECT  4.505 1.25 4.83 1.255 ;
      RECT  4.5 1.255 4.825 1.26 ;
      RECT  4.495 1.26 4.82 1.265 ;
      RECT  4.49 1.265 4.815 1.27 ;
      RECT  4.485 1.27 4.81 1.275 ;
      RECT  4.48 1.275 4.805 1.28 ;
      RECT  4.475 1.28 4.8 1.285 ;
      RECT  4.47 1.285 4.795 1.29 ;
      RECT  4.465 1.29 4.79 1.295 ;
      RECT  4.46 1.295 4.785 1.3 ;
      RECT  4.455 1.3 4.78 1.305 ;
      RECT  4.45 1.305 4.775 1.31 ;
      RECT  4.445 1.31 4.77 1.315 ;
      RECT  4.44 1.315 4.765 1.32 ;
      RECT  4.435 1.32 4.76 1.325 ;
      RECT  4.43 1.325 4.755 1.33 ;
      RECT  4.425 1.33 4.75 1.335 ;
      RECT  4.42 1.335 4.745 1.34 ;
      RECT  4.415 1.34 4.74 1.345 ;
      RECT  4.41 1.345 4.735 1.35 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.35 ;
      RECT  3.245 1.35 4.73 1.355 ;
      RECT  3.245 1.355 4.725 1.36 ;
      RECT  3.245 1.36 4.72 1.365 ;
      RECT  3.245 1.365 4.715 1.37 ;
      RECT  3.245 1.37 4.71 1.375 ;
      RECT  3.245 1.375 4.705 1.38 ;
      RECT  3.245 1.38 4.7 1.385 ;
      RECT  3.245 1.385 4.695 1.39 ;
      RECT  3.245 1.39 4.69 1.395 ;
      RECT  3.245 1.395 4.685 1.4 ;
      RECT  3.245 1.4 4.68 1.405 ;
      RECT  3.245 1.405 4.675 1.41 ;
      RECT  3.245 1.41 4.67 1.415 ;
      RECT  3.245 1.415 4.665 1.42 ;
      RECT  3.245 1.42 4.66 1.425 ;
      RECT  3.245 1.425 4.655 1.43 ;
      RECT  3.245 1.43 4.65 1.435 ;
      RECT  3.245 1.435 4.645 1.44 ;
      RECT  3.245 1.44 4.64 1.445 ;
      RECT  3.245 1.445 4.635 1.45 ;
      RECT  3.245 1.45 4.63 1.455 ;
      RECT  3.245 1.455 4.625 1.46 ;
      RECT  3.245 1.46 4.62 1.465 ;
      RECT  3.245 1.465 4.615 1.47 ;
      RECT  3.245 1.47 4.61 1.475 ;
      RECT  3.245 1.475 4.605 1.48 ;
      RECT  3.245 1.48 4.6 1.485 ;
      RECT  3.245 1.485 4.595 1.49 ;
      RECT  3.245 1.49 4.59 1.495 ;
      RECT  3.245 1.495 4.585 1.5 ;
      RECT  3.245 1.5 4.58 1.505 ;
      RECT  3.245 1.505 4.575 1.51 ;
      RECT  3.245 1.51 4.57 1.515 ;
      RECT  3.245 1.515 4.565 1.52 ;
      RECT  3.245 1.52 4.56 1.525 ;
      RECT  3.245 1.525 4.555 1.53 ;
      RECT  3.245 1.53 4.55 1.535 ;
      RECT  3.245 1.535 4.545 1.54 ;
      RECT  3.245 1.54 4.54 1.545 ;
      RECT  3.245 1.545 4.535 1.55 ;
      RECT  3.245 1.55 4.53 1.555 ;
      RECT  3.245 1.555 4.525 1.56 ;
      RECT  3.245 1.56 4.52 1.565 ;
      RECT  3.245 1.565 4.515 1.57 ;
      RECT  3.245 1.57 4.51 1.575 ;
      RECT  3.245 1.575 4.505 1.58 ;
      RECT  5.485 1.75 7.24 1.98 ;
      RECT  6.2 1.29 8.78 1.52 ;
      RECT  12.92 1.29 15.5 1.52 ;
      RECT  9.015 1.565 9.48 1.795 ;
      RECT  9.015 1.795 9.245 2.405 ;
      RECT  8.23 2.405 9.245 2.635 ;
      RECT  9.015 2.635 9.245 4.215 ;
      RECT  9.01 4.215 11.315 4.445 ;
      RECT  11.085 4.445 11.315 4.54 ;
      RECT  11.085 4.54 12.995 4.77 ;
      RECT  12.765 4.77 12.995 5.0 ;
      RECT  12.765 5.0 14.17 5.23 ;
      RECT  9.965 1.565 11.02 1.795 ;
      RECT  9.965 1.795 10.195 2.42 ;
      RECT  9.5 2.42 10.195 2.65 ;
      RECT  9.965 2.65 10.195 3.755 ;
      RECT  9.965 3.755 11.875 3.985 ;
      RECT  11.645 3.985 11.875 4.08 ;
      RECT  11.645 4.08 13.555 4.31 ;
      RECT  13.325 4.31 13.555 4.54 ;
      RECT  13.325 4.54 14.675 4.77 ;
      RECT  14.445 4.77 14.675 5.0 ;
      RECT  14.445 5.0 15.295 5.23 ;
      RECT  4.66 1.75 5.155 1.98 ;
      RECT  4.925 1.98 5.155 2.405 ;
      RECT  3.75 2.405 5.155 2.635 ;
      RECT  4.925 2.635 5.155 3.245 ;
      RECT  4.66 3.245 5.155 3.475 ;
      RECT  7.67 1.75 8.01 1.98 ;
      RECT  7.725 1.98 7.955 3.53 ;
      RECT  14.39 1.75 14.73 1.98 ;
      RECT  14.445 1.98 14.675 3.53 ;
      RECT  21.935 1.585 22.165 2.125 ;
      RECT  21.935 2.125 24.195 2.355 ;
      RECT  22.845 2.355 23.075 2.69 ;
      RECT  23.965 2.355 24.195 2.69 ;
      RECT  21.935 2.355 22.165 3.53 ;
      RECT  25.08 2.12 26.435 2.36 ;
      RECT  25.085 2.36 25.315 2.69 ;
      RECT  26.205 2.36 26.435 2.69 ;
      RECT  12.92 3.16 13.96 3.39 ;
      RECT  6.2 3.245 7.24 3.475 ;
      RECT  1.72 3.805 2.76 4.035 ;
      RECT  3.19 3.805 8.78 4.035 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  7.67 4.675 10.755 4.905 ;
      RECT  10.525 4.905 10.755 5.0 ;
      RECT  10.525 5.0 11.93 5.23 ;
      RECT  1.51 4.925 5.21 5.155 ;
      RECT  1.51 5.155 1.85 5.23 ;
      RECT  4.87 5.155 5.21 5.23 ;
  END
END MDN_FSDP_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDP_1
#      Description : D-Flip Flop w/scan, pos-edge triggered
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDP_1
  CLASS CORE ;
  FOREIGN MDN_FSDP_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 1.565 17.74 1.795 ;
      RECT  16.685 1.795 16.915 3.245 ;
      RECT  16.685 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.1 1.565 18.595 1.795 ;
      RECT  18.365 1.795 18.595 3.245 ;
      RECT  18.1 3.245 18.595 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  12.88 5.46 13.61 5.74 ;
      RECT  12.205 5.08 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 10.64 5.74 ;
      RECT  5.485 4.905 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  3.92 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.705 ;
      RECT  4.015 0.14 4.245 1.175 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.375 ;
      RECT  5.99 0.375 6.335 0.6 ;
      RECT  6.105 0.6 6.335 0.83 ;
      RECT  6.105 0.83 9.635 1.005 ;
      RECT  6.105 1.005 12.435 1.06 ;
      RECT  9.405 1.06 12.435 1.235 ;
      RECT  12.205 1.235 12.435 1.75 ;
      RECT  12.205 1.75 13.96 1.98 ;
      RECT  12.205 1.98 12.435 3.245 ;
      RECT  11.38 3.245 12.435 3.475 ;
      RECT  12.205 3.475 12.435 3.62 ;
      RECT  12.205 3.62 14.175 3.805 ;
      RECT  12.205 3.805 15.5 3.85 ;
      RECT  13.945 3.85 15.5 4.035 ;
      RECT  7.11 0.37 9.69 0.6 ;
      RECT  12.71 0.37 13.225 0.6 ;
      RECT  12.995 0.6 13.225 0.83 ;
      RECT  12.995 0.83 15.985 1.06 ;
      RECT  15.755 1.06 15.985 1.565 ;
      RECT  15.755 1.565 16.2 1.795 ;
      RECT  15.755 1.795 15.985 2.125 ;
      RECT  15.005 2.125 15.985 2.355 ;
      RECT  15.005 2.355 15.235 3.245 ;
      RECT  15.005 3.245 16.355 3.475 ;
      RECT  16.125 3.475 16.355 4.365 ;
      RECT  16.125 4.365 17.475 4.595 ;
      RECT  17.245 4.595 17.475 5.0 ;
      RECT  17.19 5.0 17.53 5.23 ;
      RECT  17.245 0.37 18.65 0.6 ;
      RECT  17.245 0.6 17.475 1.005 ;
      RECT  14.39 0.37 16.445 0.6 ;
      RECT  16.215 0.6 16.445 1.005 ;
      RECT  16.215 1.005 17.475 1.235 ;
      RECT  4.745 1.005 5.715 1.01 ;
      RECT  4.74 1.01 5.715 1.015 ;
      RECT  4.735 1.015 5.715 1.02 ;
      RECT  4.73 1.02 5.715 1.025 ;
      RECT  4.725 1.025 5.715 1.03 ;
      RECT  4.72 1.03 5.715 1.035 ;
      RECT  4.715 1.035 5.715 1.04 ;
      RECT  4.71 1.04 5.715 1.045 ;
      RECT  4.705 1.045 5.715 1.05 ;
      RECT  4.7 1.05 5.715 1.055 ;
      RECT  4.695 1.055 5.715 1.06 ;
      RECT  4.69 1.06 5.715 1.065 ;
      RECT  4.685 1.065 5.715 1.07 ;
      RECT  4.68 1.07 5.715 1.075 ;
      RECT  4.675 1.075 5.715 1.08 ;
      RECT  4.67 1.08 5.715 1.085 ;
      RECT  4.665 1.085 5.715 1.09 ;
      RECT  4.66 1.09 5.715 1.095 ;
      RECT  4.655 1.095 5.715 1.1 ;
      RECT  4.65 1.1 5.715 1.105 ;
      RECT  4.645 1.105 5.715 1.11 ;
      RECT  4.64 1.11 5.715 1.115 ;
      RECT  4.635 1.115 5.715 1.12 ;
      RECT  4.63 1.12 5.715 1.125 ;
      RECT  4.625 1.125 5.715 1.13 ;
      RECT  4.62 1.13 5.715 1.135 ;
      RECT  4.615 1.135 5.715 1.14 ;
      RECT  4.61 1.14 5.715 1.145 ;
      RECT  4.605 1.145 5.715 1.15 ;
      RECT  4.6 1.15 5.715 1.155 ;
      RECT  4.595 1.155 5.715 1.16 ;
      RECT  4.59 1.16 5.715 1.165 ;
      RECT  4.585 1.165 5.715 1.17 ;
      RECT  4.58 1.17 5.715 1.175 ;
      RECT  4.575 1.175 5.715 1.18 ;
      RECT  4.57 1.18 5.715 1.185 ;
      RECT  4.565 1.185 5.715 1.19 ;
      RECT  4.56 1.19 5.715 1.195 ;
      RECT  4.555 1.195 5.715 1.2 ;
      RECT  4.55 1.2 5.715 1.205 ;
      RECT  4.545 1.205 5.715 1.21 ;
      RECT  4.54 1.21 5.715 1.215 ;
      RECT  4.535 1.215 5.715 1.22 ;
      RECT  4.53 1.22 5.715 1.225 ;
      RECT  4.525 1.225 5.715 1.23 ;
      RECT  4.52 1.23 5.715 1.235 ;
      RECT  4.515 1.235 4.84 1.24 ;
      RECT  5.485 1.235 5.715 1.75 ;
      RECT  4.51 1.24 4.835 1.245 ;
      RECT  4.505 1.245 4.83 1.25 ;
      RECT  4.5 1.25 4.825 1.255 ;
      RECT  4.495 1.255 4.82 1.26 ;
      RECT  4.49 1.26 4.815 1.265 ;
      RECT  4.485 1.265 4.81 1.27 ;
      RECT  4.48 1.27 4.805 1.275 ;
      RECT  4.475 1.275 4.8 1.28 ;
      RECT  4.47 1.28 4.795 1.285 ;
      RECT  4.465 1.285 4.79 1.29 ;
      RECT  4.46 1.29 4.785 1.295 ;
      RECT  4.455 1.295 4.78 1.3 ;
      RECT  4.45 1.3 4.775 1.305 ;
      RECT  4.445 1.305 4.77 1.31 ;
      RECT  4.44 1.31 4.765 1.315 ;
      RECT  4.435 1.315 4.76 1.32 ;
      RECT  4.43 1.32 4.755 1.325 ;
      RECT  4.425 1.325 4.75 1.33 ;
      RECT  4.42 1.33 4.745 1.335 ;
      RECT  4.415 1.335 4.74 1.34 ;
      RECT  4.41 1.34 4.735 1.345 ;
      RECT  4.405 1.345 4.73 1.35 ;
      RECT  4.4 1.35 4.725 1.355 ;
      RECT  4.395 1.355 4.72 1.36 ;
      RECT  4.39 1.36 4.715 1.365 ;
      RECT  4.385 1.365 4.71 1.37 ;
      RECT  4.38 1.37 4.705 1.375 ;
      RECT  4.375 1.375 4.7 1.38 ;
      RECT  4.37 1.38 4.695 1.385 ;
      RECT  4.365 1.385 4.69 1.39 ;
      RECT  4.36 1.39 4.685 1.395 ;
      RECT  4.355 1.395 4.68 1.4 ;
      RECT  4.35 1.4 4.675 1.405 ;
      RECT  4.345 1.405 4.67 1.41 ;
      RECT  4.34 1.41 4.665 1.415 ;
      RECT  4.335 1.415 4.66 1.42 ;
      RECT  4.33 1.42 4.655 1.425 ;
      RECT  4.325 1.425 4.65 1.43 ;
      RECT  4.32 1.43 4.645 1.435 ;
      RECT  4.315 1.435 4.64 1.44 ;
      RECT  4.31 1.44 4.635 1.445 ;
      RECT  4.305 1.445 4.63 1.45 ;
      RECT  4.3 1.45 4.625 1.455 ;
      RECT  4.295 1.455 4.62 1.46 ;
      RECT  4.29 1.46 4.615 1.465 ;
      RECT  4.285 1.465 4.61 1.47 ;
      RECT  4.28 1.47 4.605 1.475 ;
      RECT  4.275 1.475 4.6 1.48 ;
      RECT  4.27 1.48 4.595 1.485 ;
      RECT  4.265 1.485 4.59 1.49 ;
      RECT  4.26 1.49 4.585 1.495 ;
      RECT  4.255 1.495 4.58 1.5 ;
      RECT  4.25 1.5 4.575 1.505 ;
      RECT  4.245 1.505 4.57 1.51 ;
      RECT  4.24 1.51 4.565 1.515 ;
      RECT  4.235 1.515 4.56 1.52 ;
      RECT  4.23 1.52 4.555 1.525 ;
      RECT  4.225 1.525 4.55 1.53 ;
      RECT  4.22 1.53 4.545 1.535 ;
      RECT  4.215 1.535 4.54 1.54 ;
      RECT  4.21 1.54 4.535 1.545 ;
      RECT  4.205 1.545 4.53 1.55 ;
      RECT  4.2 1.55 4.525 1.555 ;
      RECT  4.195 1.555 4.52 1.56 ;
      RECT  4.19 1.56 4.515 1.565 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  3.245 1.565 4.51 1.57 ;
      RECT  3.245 1.57 4.505 1.575 ;
      RECT  3.245 1.575 4.5 1.58 ;
      RECT  3.245 1.58 4.495 1.585 ;
      RECT  3.245 1.585 4.49 1.59 ;
      RECT  3.245 1.59 4.485 1.595 ;
      RECT  3.245 1.595 4.48 1.6 ;
      RECT  3.245 1.6 4.475 1.605 ;
      RECT  3.245 1.605 4.47 1.61 ;
      RECT  3.245 1.61 4.465 1.615 ;
      RECT  3.245 1.615 4.46 1.62 ;
      RECT  3.245 1.62 4.455 1.625 ;
      RECT  3.245 1.625 4.45 1.63 ;
      RECT  3.245 1.63 4.445 1.635 ;
      RECT  3.245 1.635 4.44 1.64 ;
      RECT  3.245 1.64 4.435 1.645 ;
      RECT  3.245 1.645 4.43 1.65 ;
      RECT  3.245 1.65 4.425 1.655 ;
      RECT  3.245 1.655 4.42 1.66 ;
      RECT  3.245 1.66 4.415 1.665 ;
      RECT  3.245 1.665 4.41 1.67 ;
      RECT  3.245 1.67 4.405 1.675 ;
      RECT  3.245 1.675 4.4 1.68 ;
      RECT  3.245 1.68 4.395 1.685 ;
      RECT  3.245 1.685 4.39 1.69 ;
      RECT  3.245 1.69 4.385 1.695 ;
      RECT  3.245 1.695 4.38 1.7 ;
      RECT  3.245 1.7 4.375 1.705 ;
      RECT  3.245 1.705 4.37 1.71 ;
      RECT  3.245 1.71 4.365 1.715 ;
      RECT  3.245 1.715 4.36 1.72 ;
      RECT  3.245 1.72 4.355 1.725 ;
      RECT  3.245 1.725 4.35 1.73 ;
      RECT  3.245 1.73 4.345 1.735 ;
      RECT  3.245 1.735 4.34 1.74 ;
      RECT  3.245 1.74 4.335 1.745 ;
      RECT  3.245 1.745 4.33 1.75 ;
      RECT  3.245 1.75 4.325 1.755 ;
      RECT  5.485 1.75 7.24 1.98 ;
      RECT  3.245 1.755 4.32 1.76 ;
      RECT  3.245 1.76 4.315 1.765 ;
      RECT  3.245 1.765 4.31 1.77 ;
      RECT  3.245 1.77 4.305 1.775 ;
      RECT  3.245 1.775 4.3 1.78 ;
      RECT  3.245 1.78 4.295 1.785 ;
      RECT  3.245 1.785 4.29 1.79 ;
      RECT  3.245 1.79 4.285 1.795 ;
      RECT  6.2 1.29 8.78 1.52 ;
      RECT  12.92 1.29 15.5 1.52 ;
      RECT  9.01 1.565 9.48 1.795 ;
      RECT  9.01 1.795 9.24 2.41 ;
      RECT  8.23 2.405 8.57 2.41 ;
      RECT  8.23 2.41 9.24 2.64 ;
      RECT  9.01 2.64 9.24 4.215 ;
      RECT  9.01 4.215 11.315 4.445 ;
      RECT  11.085 4.445 11.315 4.54 ;
      RECT  11.085 4.54 12.995 4.77 ;
      RECT  12.765 4.77 12.995 5.0 ;
      RECT  12.765 5.0 14.17 5.23 ;
      RECT  9.965 1.565 11.02 1.795 ;
      RECT  9.965 1.795 10.195 2.415 ;
      RECT  9.47 2.415 10.195 2.645 ;
      RECT  9.965 2.645 10.195 3.755 ;
      RECT  9.965 3.755 11.875 3.985 ;
      RECT  11.645 3.985 11.875 4.08 ;
      RECT  11.645 4.08 13.555 4.31 ;
      RECT  13.325 4.31 13.555 4.54 ;
      RECT  13.325 4.54 14.675 4.77 ;
      RECT  14.445 4.77 14.675 5.0 ;
      RECT  14.445 5.0 15.29 5.23 ;
      RECT  7.67 1.75 8.01 1.98 ;
      RECT  7.725 1.98 7.955 3.53 ;
      RECT  14.39 1.75 14.73 1.98 ;
      RECT  14.445 1.98 14.675 3.53 ;
      RECT  3.75 2.405 4.09 2.41 ;
      RECT  3.75 2.41 4.945 2.635 ;
      RECT  4.715 1.695 4.945 2.41 ;
      RECT  3.755 2.635 4.945 2.64 ;
      RECT  4.715 2.64 4.945 3.53 ;
      RECT  12.92 3.16 13.96 3.39 ;
      RECT  6.195 3.245 7.24 3.475 ;
      RECT  1.72 3.805 2.76 4.035 ;
      RECT  3.19 3.805 8.78 4.035 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  7.67 4.675 10.755 4.905 ;
      RECT  10.525 4.905 10.755 5.0 ;
      RECT  10.525 5.0 11.93 5.23 ;
      RECT  1.51 4.925 5.21 5.155 ;
      RECT  1.51 5.155 1.85 5.23 ;
      RECT  4.87 5.155 5.21 5.23 ;
  END
END MDN_FSDP_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDP_2
#      Description : D-Flip Flop w/scan, pos-edge triggered
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDP_2
  CLASS CORE ;
  FOREIGN MDN_FSDP_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.4 1.565 18.44 1.795 ;
      RECT  17.805 1.795 18.035 3.245 ;
      RECT  17.4 3.245 18.44 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.64 1.565 20.68 1.795 ;
      RECT  20.045 1.795 20.275 3.245 ;
      RECT  19.64 3.245 20.68 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 12.435 5.74 ;
      RECT  12.205 5.08 12.435 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.925 -0.14 20.16 0.14 ;
      RECT  18.925 0.14 19.155 0.735 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  3.92 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  4.015 0.14 4.245 1.175 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.46 0.6 ;
      RECT  6.23 0.6 6.46 0.83 ;
      RECT  6.23 0.83 9.635 1.005 ;
      RECT  6.23 1.005 12.435 1.06 ;
      RECT  9.405 1.06 12.435 1.235 ;
      RECT  12.205 1.235 12.435 1.75 ;
      RECT  12.205 1.75 13.96 1.98 ;
      RECT  12.205 1.98 12.435 3.19 ;
      RECT  11.38 3.19 12.435 3.42 ;
      RECT  12.205 3.42 12.435 3.62 ;
      RECT  12.205 3.62 14.115 3.805 ;
      RECT  12.205 3.805 15.5 3.85 ;
      RECT  13.885 3.85 15.5 4.035 ;
      RECT  7.11 0.37 9.69 0.6 ;
      RECT  12.71 0.37 13.225 0.6 ;
      RECT  12.995 0.6 13.225 0.83 ;
      RECT  12.995 0.83 15.985 1.06 ;
      RECT  15.755 1.06 15.985 1.565 ;
      RECT  15.755 1.565 16.34 1.795 ;
      RECT  16.11 1.795 16.34 2.37 ;
      RECT  16.11 2.37 17.38 2.6 ;
      RECT  16.11 2.6 16.34 3.245 ;
      RECT  15.86 3.245 16.34 3.475 ;
      RECT  17.19 0.37 18.65 0.6 ;
      RECT  19.43 0.37 20.89 0.6 ;
      RECT  19.43 0.6 19.67 1.005 ;
      RECT  14.39 0.37 16.455 0.6 ;
      RECT  16.225 0.6 16.455 1.005 ;
      RECT  16.225 1.005 19.67 1.235 ;
      RECT  4.745 1.005 5.715 1.01 ;
      RECT  4.74 1.01 5.715 1.015 ;
      RECT  4.735 1.015 5.715 1.02 ;
      RECT  4.73 1.02 5.715 1.025 ;
      RECT  4.725 1.025 5.715 1.03 ;
      RECT  4.72 1.03 5.715 1.035 ;
      RECT  4.715 1.035 5.715 1.04 ;
      RECT  4.71 1.04 5.715 1.045 ;
      RECT  4.705 1.045 5.715 1.05 ;
      RECT  4.7 1.05 5.715 1.055 ;
      RECT  4.695 1.055 5.715 1.06 ;
      RECT  4.69 1.06 5.715 1.065 ;
      RECT  4.685 1.065 5.715 1.07 ;
      RECT  4.68 1.07 5.715 1.075 ;
      RECT  4.675 1.075 5.715 1.08 ;
      RECT  4.67 1.08 5.715 1.085 ;
      RECT  4.665 1.085 5.715 1.09 ;
      RECT  4.66 1.09 5.715 1.095 ;
      RECT  4.655 1.095 5.715 1.1 ;
      RECT  4.65 1.1 5.715 1.105 ;
      RECT  4.645 1.105 5.715 1.11 ;
      RECT  4.64 1.11 5.715 1.115 ;
      RECT  4.635 1.115 5.715 1.12 ;
      RECT  4.63 1.12 5.715 1.125 ;
      RECT  4.625 1.125 5.715 1.13 ;
      RECT  4.62 1.13 5.715 1.135 ;
      RECT  4.615 1.135 5.715 1.14 ;
      RECT  4.61 1.14 5.715 1.145 ;
      RECT  4.605 1.145 5.715 1.15 ;
      RECT  4.6 1.15 5.715 1.155 ;
      RECT  4.595 1.155 5.715 1.16 ;
      RECT  4.59 1.16 5.715 1.165 ;
      RECT  4.585 1.165 5.715 1.17 ;
      RECT  4.58 1.17 5.715 1.175 ;
      RECT  4.575 1.175 5.715 1.18 ;
      RECT  4.57 1.18 5.715 1.185 ;
      RECT  4.565 1.185 5.715 1.19 ;
      RECT  4.56 1.19 5.715 1.195 ;
      RECT  4.555 1.195 5.715 1.2 ;
      RECT  4.55 1.2 5.715 1.205 ;
      RECT  4.545 1.205 5.715 1.21 ;
      RECT  4.54 1.21 5.715 1.215 ;
      RECT  4.535 1.215 5.715 1.22 ;
      RECT  4.53 1.22 5.715 1.225 ;
      RECT  4.525 1.225 5.715 1.23 ;
      RECT  4.52 1.23 5.715 1.235 ;
      RECT  4.515 1.235 4.84 1.24 ;
      RECT  5.485 1.235 5.715 1.75 ;
      RECT  4.51 1.24 4.835 1.245 ;
      RECT  4.505 1.245 4.83 1.25 ;
      RECT  4.5 1.25 4.825 1.255 ;
      RECT  4.495 1.255 4.82 1.26 ;
      RECT  4.49 1.26 4.815 1.265 ;
      RECT  4.485 1.265 4.81 1.27 ;
      RECT  4.48 1.27 4.805 1.275 ;
      RECT  4.475 1.275 4.8 1.28 ;
      RECT  4.47 1.28 4.795 1.285 ;
      RECT  4.465 1.285 4.79 1.29 ;
      RECT  4.46 1.29 4.785 1.295 ;
      RECT  4.455 1.295 4.78 1.3 ;
      RECT  4.45 1.3 4.775 1.305 ;
      RECT  4.445 1.305 4.77 1.31 ;
      RECT  4.44 1.31 4.765 1.315 ;
      RECT  4.435 1.315 4.76 1.32 ;
      RECT  4.43 1.32 4.755 1.325 ;
      RECT  4.425 1.325 4.75 1.33 ;
      RECT  4.42 1.33 4.745 1.335 ;
      RECT  4.415 1.335 4.74 1.34 ;
      RECT  4.41 1.34 4.735 1.345 ;
      RECT  4.405 1.345 4.73 1.35 ;
      RECT  4.4 1.35 4.725 1.355 ;
      RECT  4.395 1.355 4.72 1.36 ;
      RECT  4.39 1.36 4.715 1.365 ;
      RECT  4.385 1.365 4.71 1.37 ;
      RECT  4.38 1.37 4.705 1.375 ;
      RECT  4.375 1.375 4.7 1.38 ;
      RECT  4.37 1.38 4.695 1.385 ;
      RECT  4.365 1.385 4.69 1.39 ;
      RECT  4.36 1.39 4.685 1.395 ;
      RECT  4.355 1.395 4.68 1.4 ;
      RECT  4.35 1.4 4.675 1.405 ;
      RECT  4.345 1.405 4.67 1.41 ;
      RECT  4.34 1.41 4.665 1.415 ;
      RECT  4.335 1.415 4.66 1.42 ;
      RECT  4.33 1.42 4.655 1.425 ;
      RECT  4.325 1.425 4.65 1.43 ;
      RECT  4.32 1.43 4.645 1.435 ;
      RECT  4.315 1.435 4.64 1.44 ;
      RECT  4.31 1.44 4.635 1.445 ;
      RECT  4.305 1.445 4.63 1.45 ;
      RECT  4.3 1.45 4.625 1.455 ;
      RECT  4.295 1.455 4.62 1.46 ;
      RECT  4.29 1.46 4.615 1.465 ;
      RECT  4.285 1.465 4.61 1.47 ;
      RECT  4.28 1.47 4.605 1.475 ;
      RECT  4.275 1.475 4.6 1.48 ;
      RECT  4.27 1.48 4.595 1.485 ;
      RECT  4.265 1.485 4.59 1.49 ;
      RECT  4.26 1.49 4.585 1.495 ;
      RECT  4.255 1.495 4.58 1.5 ;
      RECT  4.25 1.5 4.575 1.505 ;
      RECT  4.245 1.505 4.57 1.51 ;
      RECT  4.24 1.51 4.565 1.515 ;
      RECT  4.235 1.515 4.56 1.52 ;
      RECT  4.23 1.52 4.555 1.525 ;
      RECT  4.225 1.525 4.55 1.53 ;
      RECT  4.22 1.53 4.545 1.535 ;
      RECT  4.215 1.535 4.54 1.54 ;
      RECT  4.21 1.54 4.535 1.545 ;
      RECT  4.205 1.545 4.53 1.55 ;
      RECT  4.2 1.55 4.525 1.555 ;
      RECT  4.195 1.555 4.52 1.56 ;
      RECT  4.19 1.56 4.515 1.565 ;
      RECT  4.185 1.565 4.51 1.57 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.57 ;
      RECT  3.245 1.57 4.505 1.575 ;
      RECT  3.245 1.575 4.5 1.58 ;
      RECT  3.245 1.58 4.495 1.585 ;
      RECT  3.245 1.585 4.49 1.59 ;
      RECT  3.245 1.59 4.485 1.595 ;
      RECT  3.245 1.595 4.48 1.6 ;
      RECT  3.245 1.6 4.475 1.605 ;
      RECT  3.245 1.605 4.47 1.61 ;
      RECT  3.245 1.61 4.465 1.615 ;
      RECT  3.245 1.615 4.46 1.62 ;
      RECT  3.245 1.62 4.455 1.625 ;
      RECT  3.245 1.625 4.45 1.63 ;
      RECT  3.245 1.63 4.445 1.635 ;
      RECT  3.245 1.635 4.44 1.64 ;
      RECT  3.245 1.64 4.435 1.645 ;
      RECT  3.245 1.645 4.43 1.65 ;
      RECT  3.245 1.65 4.425 1.655 ;
      RECT  3.245 1.655 4.42 1.66 ;
      RECT  3.245 1.66 4.415 1.665 ;
      RECT  3.245 1.665 4.41 1.67 ;
      RECT  3.245 1.67 4.405 1.675 ;
      RECT  3.245 1.675 4.4 1.68 ;
      RECT  3.245 1.68 4.395 1.685 ;
      RECT  3.245 1.685 4.39 1.69 ;
      RECT  3.245 1.69 4.385 1.695 ;
      RECT  3.245 1.695 4.38 1.7 ;
      RECT  3.245 1.7 4.375 1.705 ;
      RECT  3.245 1.705 4.37 1.71 ;
      RECT  3.245 1.71 4.365 1.715 ;
      RECT  3.245 1.715 4.36 1.72 ;
      RECT  3.245 1.72 4.355 1.725 ;
      RECT  3.245 1.725 4.35 1.73 ;
      RECT  3.245 1.73 4.345 1.735 ;
      RECT  3.245 1.735 4.34 1.74 ;
      RECT  3.245 1.74 4.335 1.745 ;
      RECT  3.245 1.745 4.33 1.75 ;
      RECT  3.245 1.75 4.325 1.755 ;
      RECT  5.485 1.75 7.24 1.98 ;
      RECT  3.245 1.755 4.32 1.76 ;
      RECT  3.245 1.76 4.315 1.765 ;
      RECT  3.245 1.765 4.31 1.77 ;
      RECT  3.245 1.77 4.305 1.775 ;
      RECT  3.245 1.775 4.3 1.78 ;
      RECT  3.245 1.78 4.295 1.785 ;
      RECT  3.245 1.785 4.29 1.79 ;
      RECT  3.245 1.79 4.285 1.795 ;
      RECT  3.245 1.795 4.28 1.8 ;
      RECT  6.2 1.29 8.78 1.52 ;
      RECT  12.92 1.29 15.5 1.52 ;
      RECT  9.01 1.565 9.48 1.795 ;
      RECT  9.01 1.795 9.24 2.395 ;
      RECT  8.23 2.395 9.24 2.625 ;
      RECT  9.01 2.625 9.24 4.215 ;
      RECT  9.01 4.215 11.315 4.445 ;
      RECT  11.085 4.445 11.315 4.54 ;
      RECT  11.085 4.54 12.995 4.77 ;
      RECT  12.765 4.77 12.995 5.0 ;
      RECT  12.765 5.0 14.17 5.23 ;
      RECT  9.965 1.565 11.02 1.795 ;
      RECT  9.965 1.795 10.195 2.415 ;
      RECT  9.475 2.415 10.195 2.645 ;
      RECT  9.965 2.645 10.195 3.755 ;
      RECT  9.965 3.755 11.875 3.985 ;
      RECT  11.645 3.985 11.875 4.08 ;
      RECT  11.645 4.08 13.555 4.31 ;
      RECT  13.325 4.31 13.555 4.365 ;
      RECT  13.325 4.365 14.675 4.595 ;
      RECT  14.445 4.595 14.675 5.0 ;
      RECT  14.445 5.0 15.29 5.23 ;
      RECT  7.665 1.75 8.005 1.98 ;
      RECT  7.725 1.98 7.955 3.53 ;
      RECT  14.39 1.75 14.73 1.98 ;
      RECT  14.445 1.98 14.675 3.53 ;
      RECT  4.715 1.695 4.945 2.41 ;
      RECT  3.75 2.41 4.945 2.64 ;
      RECT  4.715 2.64 4.945 3.53 ;
      RECT  12.92 3.16 13.96 3.39 ;
      RECT  6.2 3.245 7.24 3.475 ;
      RECT  1.72 3.805 2.76 4.035 ;
      RECT  3.19 3.805 8.78 4.035 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  7.67 4.675 10.755 4.905 ;
      RECT  10.525 4.905 10.755 5.0 ;
      RECT  10.525 5.0 11.93 5.23 ;
      RECT  1.51 4.925 5.21 5.155 ;
      RECT  1.51 5.155 1.85 5.23 ;
      RECT  4.87 5.155 5.21 5.23 ;
  END
END MDN_FSDP_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDPHRBQ_1
#      Description : D-Flip Flop w/scan, pos-edge triggered, lo-async-clear, sync hold, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(iq&EN&!SE)|(!EN&(!SE&D))|(SE&SI),clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDPHRBQ_1
  CLASS CORE ;
  FOREIGN MDN_FSDPHRBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 26.88 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  26.18 2.125 26.46 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 8.54 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 11.9 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  24.12 1.565 24.755 1.795 ;
      RECT  24.525 1.795 24.755 3.245 ;
      RECT  24.12 3.245 24.755 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.22 2.125 18.62 2.355 ;
      RECT  17.22 2.355 17.5 2.915 ;
      RECT  18.34 2.355 18.62 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 4.87 25.875 5.46 ;
      RECT  25.645 5.46 27.05 5.74 ;
      RECT  23.405 4.87 23.635 5.46 ;
      RECT  22.96 5.46 23.635 5.74 ;
      RECT  18.925 5.0 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  16.685 5.08 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 26.88 5.74 ;
      LAYER VIA12 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 -0.14 27.05 0.14 ;
      RECT  25.645 0.14 25.875 0.73 ;
      RECT  23.405 -0.14 24.08 0.14 ;
      RECT  23.405 0.14 23.635 0.6 ;
      RECT  17.36 -0.14 18.48 0.14 ;
      RECT  17.805 0.14 18.035 1.005 ;
      RECT  17.4 1.005 18.44 1.235 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 26.88 0.14 ;
      LAYER VIA12 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  18.07 -0.13 18.33 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  7.11 0.37 7.45 0.445 ;
      RECT  7.11 0.445 11.61 0.675 ;
      RECT  11.38 0.675 11.61 1.005 ;
      RECT  11.38 1.005 12.435 1.235 ;
      RECT  12.205 1.235 12.435 3.245 ;
      RECT  11.38 3.245 12.435 3.475 ;
      RECT  20.55 0.37 20.89 0.83 ;
      RECT  18.67 0.83 24.195 1.005 ;
      RECT  18.67 1.005 25.315 1.06 ;
      RECT  23.965 1.06 25.315 1.235 ;
      RECT  18.67 1.06 18.9 1.565 ;
      RECT  25.085 1.235 25.315 3.805 ;
      RECT  13.83 0.37 17.12 0.6 ;
      RECT  16.89 0.6 17.12 1.565 ;
      RECT  16.89 1.565 18.9 1.795 ;
      RECT  24.82 3.805 25.315 4.035 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 1.565 ;
      RECT  1.005 1.565 2.76 1.795 ;
      RECT  1.72 1.005 4.035 1.235 ;
      RECT  3.805 1.235 4.035 2.125 ;
      RECT  3.805 2.125 6.275 2.355 ;
      RECT  6.045 2.355 6.275 2.69 ;
      RECT  3.805 2.355 4.035 3.805 ;
      RECT  1.72 3.805 4.035 4.035 ;
      RECT  6.2 1.005 11.02 1.235 ;
      RECT  25.645 1.005 26.7 1.235 ;
      RECT  25.645 1.235 25.875 4.365 ;
      RECT  23.965 4.365 26.7 4.41 ;
      RECT  20.605 4.41 26.7 4.54 ;
      RECT  16.565 4.54 26.7 4.545 ;
      RECT  16.56 4.545 26.7 4.55 ;
      RECT  16.555 4.55 26.7 4.555 ;
      RECT  16.55 4.555 26.7 4.56 ;
      RECT  16.545 4.56 26.7 4.565 ;
      RECT  16.54 4.565 26.7 4.57 ;
      RECT  16.535 4.57 26.7 4.575 ;
      RECT  16.53 4.575 26.7 4.58 ;
      RECT  16.525 4.58 26.7 4.585 ;
      RECT  16.52 4.585 26.7 4.59 ;
      RECT  16.515 4.59 26.7 4.595 ;
      RECT  16.51 4.595 24.195 4.6 ;
      RECT  25.03 4.595 25.26 5.0 ;
      RECT  16.505 4.6 24.195 4.605 ;
      RECT  16.5 4.605 24.195 4.61 ;
      RECT  16.495 4.61 24.195 4.615 ;
      RECT  16.49 4.615 24.195 4.62 ;
      RECT  16.485 4.62 24.195 4.625 ;
      RECT  16.48 4.625 24.195 4.63 ;
      RECT  16.475 4.63 24.195 4.635 ;
      RECT  16.47 4.635 24.195 4.64 ;
      RECT  16.465 4.64 20.835 4.645 ;
      RECT  21.68 4.64 21.91 5.0 ;
      RECT  16.46 4.645 20.835 4.65 ;
      RECT  16.455 4.65 20.835 4.655 ;
      RECT  16.45 4.655 20.835 4.66 ;
      RECT  16.445 4.66 20.835 4.665 ;
      RECT  16.44 4.665 20.835 4.67 ;
      RECT  16.435 4.67 20.835 4.675 ;
      RECT  16.43 4.675 20.835 4.68 ;
      RECT  16.425 4.68 20.835 4.685 ;
      RECT  16.42 4.685 20.835 4.69 ;
      RECT  16.415 4.69 20.835 4.695 ;
      RECT  16.41 4.695 20.835 4.7 ;
      RECT  16.405 4.7 20.835 4.705 ;
      RECT  16.4 4.705 20.835 4.71 ;
      RECT  16.395 4.71 20.835 4.715 ;
      RECT  16.39 4.715 20.835 4.72 ;
      RECT  16.385 4.72 20.835 4.725 ;
      RECT  16.38 4.725 20.835 4.73 ;
      RECT  16.375 4.73 20.835 4.735 ;
      RECT  16.37 4.735 20.835 4.74 ;
      RECT  16.365 4.74 20.835 4.745 ;
      RECT  16.36 4.745 20.835 4.75 ;
      RECT  16.355 4.75 20.835 4.755 ;
      RECT  16.35 4.755 20.835 4.76 ;
      RECT  16.345 4.76 20.835 4.765 ;
      RECT  16.34 4.765 20.835 4.77 ;
      RECT  16.335 4.77 16.66 4.775 ;
      RECT  16.33 4.775 16.655 4.78 ;
      RECT  16.325 4.78 16.65 4.785 ;
      RECT  16.32 4.785 16.645 4.79 ;
      RECT  16.315 4.79 16.64 4.795 ;
      RECT  16.31 4.795 16.635 4.8 ;
      RECT  16.305 4.8 16.63 4.805 ;
      RECT  16.3 4.805 16.625 4.81 ;
      RECT  16.295 4.81 16.62 4.815 ;
      RECT  16.29 4.815 16.615 4.82 ;
      RECT  16.285 4.82 16.61 4.825 ;
      RECT  16.28 4.825 16.605 4.83 ;
      RECT  16.275 4.83 16.6 4.835 ;
      RECT  16.27 4.835 16.595 4.84 ;
      RECT  16.265 4.84 16.59 4.845 ;
      RECT  16.26 4.845 16.585 4.85 ;
      RECT  16.255 4.85 16.58 4.855 ;
      RECT  16.25 4.855 16.575 4.86 ;
      RECT  16.245 4.86 16.57 4.865 ;
      RECT  16.24 4.865 16.565 4.87 ;
      RECT  16.235 4.87 16.56 4.875 ;
      RECT  16.23 4.875 16.555 4.88 ;
      RECT  16.225 4.88 16.55 4.885 ;
      RECT  16.22 4.885 16.545 4.89 ;
      RECT  16.215 4.89 16.54 4.895 ;
      RECT  16.21 4.895 16.535 4.9 ;
      RECT  16.205 4.9 16.53 4.905 ;
      RECT  16.2 4.905 16.525 4.91 ;
      RECT  16.195 4.91 16.52 4.915 ;
      RECT  16.19 4.915 16.515 4.92 ;
      RECT  16.185 4.92 16.51 4.925 ;
      RECT  16.18 4.925 16.505 4.93 ;
      RECT  16.175 4.93 16.5 4.935 ;
      RECT  16.17 4.935 16.495 4.94 ;
      RECT  16.165 4.94 16.49 4.945 ;
      RECT  16.16 4.945 16.485 4.95 ;
      RECT  16.155 4.95 16.48 4.955 ;
      RECT  16.15 4.955 16.475 4.96 ;
      RECT  16.145 4.96 16.47 4.965 ;
      RECT  16.14 4.965 16.465 4.97 ;
      RECT  16.135 4.97 16.46 4.975 ;
      RECT  16.13 4.975 16.455 4.98 ;
      RECT  16.125 4.98 16.45 4.985 ;
      RECT  16.12 4.985 16.445 4.99 ;
      RECT  16.115 4.99 16.44 4.995 ;
      RECT  16.11 4.995 16.435 5.0 ;
      RECT  14.96 5.0 16.43 5.005 ;
      RECT  21.68 5.0 22.02 5.23 ;
      RECT  25.03 5.0 25.37 5.23 ;
      RECT  14.96 5.005 16.425 5.01 ;
      RECT  14.96 5.01 16.42 5.015 ;
      RECT  14.96 5.015 16.415 5.02 ;
      RECT  14.96 5.02 16.41 5.025 ;
      RECT  14.96 5.025 16.405 5.03 ;
      RECT  14.96 5.03 16.4 5.035 ;
      RECT  14.96 5.035 16.395 5.04 ;
      RECT  14.96 5.04 16.39 5.045 ;
      RECT  14.96 5.045 16.385 5.05 ;
      RECT  14.96 5.05 16.38 5.055 ;
      RECT  14.96 5.055 16.375 5.06 ;
      RECT  14.96 5.06 16.37 5.065 ;
      RECT  14.96 5.065 16.365 5.07 ;
      RECT  14.96 5.07 16.36 5.075 ;
      RECT  14.96 5.075 16.355 5.08 ;
      RECT  14.96 5.08 16.35 5.085 ;
      RECT  14.96 5.085 16.345 5.09 ;
      RECT  14.96 5.09 16.34 5.095 ;
      RECT  14.96 5.095 16.335 5.1 ;
      RECT  14.96 5.1 16.33 5.105 ;
      RECT  14.96 5.105 16.325 5.11 ;
      RECT  14.96 5.11 16.32 5.115 ;
      RECT  14.96 5.115 16.315 5.12 ;
      RECT  14.96 5.12 16.31 5.125 ;
      RECT  14.96 5.125 16.305 5.13 ;
      RECT  14.96 5.13 16.3 5.135 ;
      RECT  14.96 5.135 16.295 5.14 ;
      RECT  14.96 5.14 16.29 5.145 ;
      RECT  14.96 5.145 16.285 5.15 ;
      RECT  14.96 5.15 16.28 5.155 ;
      RECT  14.96 5.155 16.275 5.16 ;
      RECT  14.96 5.16 16.27 5.165 ;
      RECT  14.96 5.165 16.265 5.17 ;
      RECT  14.96 5.17 16.26 5.175 ;
      RECT  14.96 5.175 16.255 5.18 ;
      RECT  14.96 5.18 16.25 5.185 ;
      RECT  14.96 5.185 16.245 5.19 ;
      RECT  14.96 5.19 16.24 5.195 ;
      RECT  14.96 5.195 16.235 5.2 ;
      RECT  14.96 5.2 16.23 5.205 ;
      RECT  14.96 5.205 16.225 5.21 ;
      RECT  14.96 5.21 16.22 5.215 ;
      RECT  14.96 5.215 16.215 5.22 ;
      RECT  14.96 5.22 16.21 5.225 ;
      RECT  14.96 5.225 16.205 5.23 ;
      RECT  13.62 1.29 16.2 1.52 ;
      RECT  19.64 1.29 23.635 1.52 ;
      RECT  23.405 1.52 23.635 2.405 ;
      RECT  23.015 2.405 24.16 2.635 ;
      RECT  23.405 2.635 23.635 3.95 ;
      RECT  20.16 3.95 23.635 4.065 ;
      RECT  18.1 4.065 23.635 4.18 ;
      RECT  18.1 4.18 20.39 4.295 ;
      RECT  14.39 1.75 14.73 1.98 ;
      RECT  14.39 1.98 14.62 2.975 ;
      RECT  14.39 2.975 14.675 3.315 ;
      RECT  15.005 1.75 15.5 1.98 ;
      RECT  15.005 1.98 15.235 3.15 ;
      RECT  14.905 3.15 15.235 3.375 ;
      RECT  14.905 3.375 15.135 3.56 ;
      RECT  13.73 3.56 15.135 3.79 ;
      RECT  13.73 3.79 13.96 3.805 ;
      RECT  3.19 0.445 4.595 0.675 ;
      RECT  4.365 0.675 4.595 1.565 ;
      RECT  4.365 1.565 9.48 1.795 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  7.67 3.245 10.195 3.475 ;
      RECT  9.965 3.475 10.195 3.805 ;
      RECT  9.965 3.805 13.96 4.035 ;
      RECT  19.13 1.75 20.68 1.98 ;
      RECT  19.13 1.98 19.36 3.03 ;
      RECT  18.925 3.03 22.22 3.145 ;
      RECT  12.765 0.83 16.66 1.06 ;
      RECT  12.765 1.06 12.995 1.565 ;
      RECT  16.43 1.06 16.66 2.405 ;
      RECT  12.765 1.565 13.26 1.795 ;
      RECT  12.765 1.795 12.995 3.245 ;
      RECT  16.07 2.405 16.66 2.635 ;
      RECT  16.43 2.635 16.66 3.145 ;
      RECT  16.43 3.145 22.22 3.26 ;
      RECT  12.765 3.245 13.26 3.475 ;
      RECT  16.43 3.26 19.155 3.375 ;
      RECT  21.11 1.75 21.45 1.98 ;
      RECT  21.11 1.98 21.34 2.405 ;
      RECT  19.59 2.405 21.34 2.635 ;
      RECT  21.88 1.75 22.92 1.98 ;
      RECT  22.45 1.98 22.68 3.49 ;
      RECT  19.62 3.49 22.92 3.605 ;
      RECT  15.365 3.605 22.92 3.72 ;
      RECT  15.365 3.72 19.88 3.835 ;
      RECT  15.365 3.835 15.595 4.02 ;
      RECT  14.445 4.02 15.595 4.25 ;
      RECT  14.445 4.25 14.675 4.365 ;
      RECT  11.745 4.365 14.675 4.595 ;
      RECT  11.745 4.595 11.975 5.0 ;
      RECT  10.48 5.0 11.975 5.23 ;
      RECT  3.245 1.51 3.475 3.53 ;
      RECT  8.44 3.805 9.48 4.035 ;
      RECT  15.825 4.065 17.74 4.295 ;
      RECT  15.825 4.295 16.055 4.48 ;
      RECT  15.16 4.48 16.055 4.71 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.66 4.365 6.275 4.595 ;
      RECT  6.045 4.595 6.275 4.985 ;
      RECT  6.045 4.985 10.25 5.215 ;
      RECT  6.9 4.365 11.02 4.595 ;
      RECT  1.51 5.0 5.21 5.23 ;
      RECT  12.71 5.0 14.73 5.23 ;
      RECT  19.43 5.0 21.45 5.23 ;
  END
END MDN_FSDPHRBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDPHRBQ_2
#      Description : D-Flip Flop w/scan, pos-edge triggered, lo-async-clear, sync hold, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(iq&EN&!SE)|(!EN&(!SE&D))|(SE&SI),clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDPHRBQ_2
  CLASS CORE ;
  FOREIGN MDN_FSDPHRBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 29.12 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  27.27 0.37 27.61 0.6 ;
      RECT  27.3 0.6 27.58 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 2.1 8.515 2.38 ;
      RECT  8.285 2.38 8.515 2.69 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 11.9 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  24.12 1.565 25.16 1.795 ;
      RECT  24.525 1.795 24.755 3.245 ;
      RECT  24.12 3.245 25.16 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.22 2.125 18.62 2.355 ;
      RECT  17.22 2.355 17.5 2.915 ;
      RECT  18.34 2.355 18.62 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 2.94 2.355 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  27.885 4.9 28.115 5.46 ;
      RECT  27.885 5.46 29.29 5.74 ;
      RECT  25.645 4.87 25.875 5.46 ;
      RECT  25.645 5.46 26.32 5.74 ;
      RECT  23.405 4.87 23.635 5.46 ;
      RECT  22.96 5.46 23.635 5.74 ;
      RECT  18.925 5.08 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 5.08 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 29.12 5.74 ;
      LAYER VIA12 ;
      RECT  28.15 5.47 28.41 5.73 ;
      RECT  28.71 5.47 28.97 5.73 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  27.885 -0.14 29.29 0.14 ;
      RECT  27.885 0.14 28.115 0.7 ;
      RECT  23.405 -0.14 25.875 0.14 ;
      RECT  23.405 0.14 23.635 0.6 ;
      RECT  25.645 0.14 25.875 0.73 ;
      RECT  17.36 -0.14 18.09 0.14 ;
      RECT  17.805 0.14 18.035 1.005 ;
      RECT  17.4 1.005 18.44 1.235 ;
      RECT  11.03 -0.14 12.435 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 29.12 0.14 ;
      LAYER VIA12 ;
      RECT  28.15 -0.13 28.41 0.13 ;
      RECT  28.71 -0.13 28.97 0.13 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  24.79 -0.13 25.05 0.13 ;
      RECT  25.35 -0.13 25.61 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  7.11 0.37 7.45 0.445 ;
      RECT  7.11 0.445 11.61 0.675 ;
      RECT  11.38 0.675 11.61 1.005 ;
      RECT  11.38 1.005 12.435 1.235 ;
      RECT  12.205 1.235 12.435 3.245 ;
      RECT  11.38 3.245 12.435 3.475 ;
      RECT  23.91 0.37 25.37 0.6 ;
      RECT  3.19 0.445 4.595 0.675 ;
      RECT  4.365 0.675 4.595 1.565 ;
      RECT  4.365 1.565 9.48 1.795 ;
      RECT  8.845 1.795 9.075 3.03 ;
      RECT  7.67 3.03 9.075 3.26 ;
      RECT  20.55 0.37 20.89 0.83 ;
      RECT  18.67 0.83 24.195 1.005 ;
      RECT  18.67 1.005 25.875 1.06 ;
      RECT  23.965 1.06 25.875 1.235 ;
      RECT  18.67 1.06 18.9 1.565 ;
      RECT  25.645 1.235 25.875 1.565 ;
      RECT  13.83 0.37 17.12 0.6 ;
      RECT  16.89 0.6 17.12 1.565 ;
      RECT  16.89 1.565 18.9 1.795 ;
      RECT  25.645 1.565 26.7 1.795 ;
      RECT  25.645 1.795 25.875 3.245 ;
      RECT  25.645 3.245 26.7 3.475 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 1.565 ;
      RECT  1.005 1.565 2.76 1.795 ;
      RECT  1.72 1.005 4.035 1.235 ;
      RECT  3.805 1.235 4.035 2.125 ;
      RECT  3.805 2.125 6.275 2.355 ;
      RECT  6.045 2.355 6.275 2.69 ;
      RECT  3.805 2.355 4.035 3.805 ;
      RECT  1.72 3.805 4.035 4.035 ;
      RECT  6.2 1.005 11.02 1.235 ;
      RECT  13.62 1.29 16.2 1.52 ;
      RECT  19.64 1.29 23.635 1.52 ;
      RECT  23.405 1.52 23.635 2.405 ;
      RECT  22.99 2.405 24.175 2.635 ;
      RECT  23.405 2.635 23.635 3.95 ;
      RECT  20.045 3.95 23.635 4.065 ;
      RECT  18.1 4.065 23.635 4.18 ;
      RECT  18.1 4.18 20.275 4.295 ;
      RECT  27.06 1.565 27.555 1.795 ;
      RECT  27.325 1.795 27.555 2.405 ;
      RECT  26.15 2.405 27.555 2.635 ;
      RECT  27.325 2.635 27.555 3.245 ;
      RECT  27.06 3.245 27.555 3.475 ;
      RECT  14.39 1.75 14.73 1.98 ;
      RECT  14.39 1.98 14.62 2.99 ;
      RECT  14.39 2.99 14.675 3.33 ;
      RECT  15.005 1.75 15.5 1.98 ;
      RECT  15.005 1.98 15.235 3.19 ;
      RECT  14.915 3.19 15.235 3.42 ;
      RECT  14.915 3.42 15.145 3.56 ;
      RECT  13.885 3.56 15.145 3.79 ;
      RECT  13.885 3.79 14.115 3.805 ;
      RECT  9.965 3.805 14.115 3.95 ;
      RECT  7.67 3.95 14.115 4.035 ;
      RECT  7.67 4.035 10.195 4.18 ;
      RECT  19.13 1.75 20.68 1.98 ;
      RECT  19.13 1.98 19.36 3.03 ;
      RECT  18.925 3.03 22.22 3.145 ;
      RECT  12.765 0.83 16.66 1.06 ;
      RECT  12.765 1.06 12.995 1.565 ;
      RECT  16.43 1.06 16.66 2.405 ;
      RECT  12.765 1.565 13.26 1.795 ;
      RECT  12.765 1.795 12.995 3.245 ;
      RECT  16.07 2.405 16.66 2.635 ;
      RECT  16.43 2.635 16.66 3.145 ;
      RECT  16.43 3.145 22.22 3.26 ;
      RECT  12.765 3.245 13.26 3.475 ;
      RECT  16.43 3.26 19.155 3.375 ;
      RECT  21.11 1.75 21.45 1.98 ;
      RECT  21.11 1.98 21.34 2.405 ;
      RECT  19.59 2.405 21.34 2.635 ;
      RECT  21.88 1.75 22.92 1.98 ;
      RECT  22.53 1.98 22.76 3.49 ;
      RECT  19.485 3.49 22.92 3.605 ;
      RECT  15.375 3.605 22.92 3.72 ;
      RECT  15.375 3.72 19.715 3.835 ;
      RECT  15.375 3.835 15.605 4.02 ;
      RECT  14.445 4.02 15.605 4.25 ;
      RECT  14.445 4.25 14.675 4.365 ;
      RECT  11.645 4.365 14.675 4.595 ;
      RECT  11.645 4.595 11.875 5.0 ;
      RECT  10.48 5.0 11.875 5.215 ;
      RECT  10.48 5.215 11.87 5.23 ;
      RECT  3.245 1.51 3.475 3.53 ;
      RECT  8.44 3.49 9.48 3.72 ;
      RECT  15.835 4.07 17.74 4.3 ;
      RECT  15.835 4.3 16.065 4.48 ;
      RECT  15.16 4.48 16.065 4.71 ;
      RECT  20.6 4.41 26.38 4.54 ;
      RECT  16.565 4.54 26.38 4.545 ;
      RECT  16.56 4.545 26.38 4.55 ;
      RECT  16.555 4.55 26.38 4.555 ;
      RECT  16.55 4.555 26.38 4.56 ;
      RECT  16.545 4.56 26.38 4.565 ;
      RECT  16.54 4.565 26.38 4.57 ;
      RECT  16.535 4.57 26.38 4.575 ;
      RECT  16.53 4.575 26.38 4.58 ;
      RECT  16.525 4.58 26.38 4.585 ;
      RECT  16.52 4.585 26.38 4.59 ;
      RECT  16.515 4.59 26.38 4.595 ;
      RECT  16.51 4.595 26.38 4.6 ;
      RECT  16.505 4.6 26.38 4.605 ;
      RECT  16.5 4.605 26.38 4.61 ;
      RECT  16.495 4.61 26.38 4.615 ;
      RECT  16.49 4.615 26.38 4.62 ;
      RECT  16.485 4.62 26.38 4.625 ;
      RECT  16.48 4.625 26.38 4.63 ;
      RECT  16.475 4.63 26.38 4.635 ;
      RECT  16.47 4.635 26.38 4.64 ;
      RECT  16.465 4.64 20.845 4.645 ;
      RECT  21.68 4.64 21.91 5.0 ;
      RECT  26.15 4.64 26.38 5.0 ;
      RECT  16.46 4.645 20.845 4.65 ;
      RECT  16.455 4.65 20.845 4.655 ;
      RECT  16.45 4.655 20.845 4.66 ;
      RECT  16.445 4.66 20.845 4.665 ;
      RECT  16.44 4.665 20.845 4.67 ;
      RECT  16.435 4.67 20.845 4.675 ;
      RECT  16.43 4.675 20.845 4.68 ;
      RECT  16.425 4.68 20.845 4.685 ;
      RECT  16.42 4.685 20.845 4.69 ;
      RECT  16.415 4.69 20.845 4.695 ;
      RECT  16.41 4.695 20.845 4.7 ;
      RECT  16.405 4.7 20.845 4.705 ;
      RECT  16.4 4.705 20.845 4.71 ;
      RECT  16.395 4.71 20.845 4.715 ;
      RECT  16.39 4.715 20.845 4.72 ;
      RECT  16.385 4.72 20.845 4.725 ;
      RECT  16.38 4.725 20.845 4.73 ;
      RECT  16.375 4.73 20.845 4.735 ;
      RECT  16.37 4.735 20.845 4.74 ;
      RECT  16.365 4.74 20.845 4.745 ;
      RECT  16.36 4.745 20.845 4.75 ;
      RECT  16.355 4.75 20.845 4.755 ;
      RECT  16.35 4.755 20.845 4.76 ;
      RECT  16.345 4.76 20.845 4.765 ;
      RECT  16.34 4.765 20.845 4.77 ;
      RECT  16.335 4.77 16.66 4.775 ;
      RECT  16.33 4.775 16.655 4.78 ;
      RECT  16.325 4.78 16.65 4.785 ;
      RECT  16.32 4.785 16.645 4.79 ;
      RECT  16.315 4.79 16.64 4.795 ;
      RECT  16.31 4.795 16.635 4.8 ;
      RECT  16.305 4.8 16.63 4.805 ;
      RECT  16.3 4.805 16.625 4.81 ;
      RECT  16.295 4.81 16.62 4.815 ;
      RECT  16.29 4.815 16.615 4.82 ;
      RECT  16.285 4.82 16.61 4.825 ;
      RECT  16.28 4.825 16.605 4.83 ;
      RECT  16.275 4.83 16.6 4.835 ;
      RECT  16.27 4.835 16.595 4.84 ;
      RECT  16.265 4.84 16.59 4.845 ;
      RECT  16.26 4.845 16.585 4.85 ;
      RECT  16.255 4.85 16.58 4.855 ;
      RECT  16.25 4.855 16.575 4.86 ;
      RECT  16.245 4.86 16.57 4.865 ;
      RECT  16.24 4.865 16.565 4.87 ;
      RECT  16.235 4.87 16.56 4.875 ;
      RECT  16.23 4.875 16.555 4.88 ;
      RECT  16.225 4.88 16.55 4.885 ;
      RECT  16.22 4.885 16.545 4.89 ;
      RECT  16.215 4.89 16.54 4.895 ;
      RECT  16.21 4.895 16.535 4.9 ;
      RECT  16.205 4.9 16.53 4.905 ;
      RECT  16.2 4.905 16.525 4.91 ;
      RECT  16.195 4.91 16.52 4.915 ;
      RECT  16.19 4.915 16.515 4.92 ;
      RECT  16.185 4.92 16.51 4.925 ;
      RECT  16.18 4.925 16.505 4.93 ;
      RECT  16.175 4.93 16.5 4.935 ;
      RECT  16.17 4.935 16.495 4.94 ;
      RECT  16.165 4.94 16.49 4.945 ;
      RECT  16.16 4.945 16.485 4.95 ;
      RECT  16.155 4.95 16.48 4.955 ;
      RECT  16.15 4.955 16.475 4.96 ;
      RECT  16.145 4.96 16.47 4.965 ;
      RECT  16.14 4.965 16.465 4.97 ;
      RECT  16.135 4.97 16.46 4.975 ;
      RECT  16.13 4.975 16.455 4.98 ;
      RECT  16.125 4.98 16.45 4.985 ;
      RECT  16.12 4.985 16.445 4.99 ;
      RECT  16.115 4.99 16.44 4.995 ;
      RECT  16.11 4.995 16.435 5.0 ;
      RECT  14.95 5.0 16.43 5.005 ;
      RECT  21.68 5.0 22.02 5.23 ;
      RECT  26.15 5.0 26.49 5.23 ;
      RECT  14.95 5.005 16.425 5.01 ;
      RECT  14.95 5.01 16.42 5.015 ;
      RECT  14.95 5.015 16.415 5.02 ;
      RECT  14.95 5.02 16.41 5.025 ;
      RECT  14.95 5.025 16.405 5.03 ;
      RECT  14.95 5.03 16.4 5.035 ;
      RECT  14.95 5.035 16.395 5.04 ;
      RECT  14.95 5.04 16.39 5.045 ;
      RECT  14.95 5.045 16.385 5.05 ;
      RECT  14.95 5.05 16.38 5.055 ;
      RECT  14.95 5.055 16.375 5.06 ;
      RECT  14.95 5.06 16.37 5.065 ;
      RECT  14.95 5.065 16.365 5.07 ;
      RECT  14.95 5.07 16.36 5.075 ;
      RECT  14.95 5.075 16.355 5.08 ;
      RECT  14.95 5.08 16.35 5.085 ;
      RECT  14.95 5.085 16.345 5.09 ;
      RECT  14.95 5.09 16.34 5.095 ;
      RECT  14.95 5.095 16.335 5.1 ;
      RECT  14.95 5.1 16.33 5.105 ;
      RECT  14.95 5.105 16.325 5.11 ;
      RECT  14.95 5.11 16.32 5.115 ;
      RECT  14.95 5.115 16.315 5.12 ;
      RECT  14.95 5.12 16.31 5.125 ;
      RECT  14.95 5.125 16.305 5.13 ;
      RECT  14.95 5.13 16.3 5.135 ;
      RECT  14.95 5.135 16.295 5.14 ;
      RECT  14.95 5.14 16.29 5.145 ;
      RECT  14.95 5.145 16.285 5.15 ;
      RECT  14.95 5.15 16.28 5.155 ;
      RECT  14.95 5.155 16.275 5.16 ;
      RECT  14.95 5.16 16.27 5.165 ;
      RECT  14.95 5.165 16.265 5.17 ;
      RECT  14.95 5.17 16.26 5.175 ;
      RECT  14.95 5.175 16.255 5.18 ;
      RECT  14.95 5.18 16.25 5.185 ;
      RECT  14.95 5.185 16.245 5.19 ;
      RECT  14.95 5.19 16.24 5.195 ;
      RECT  14.95 5.195 16.235 5.2 ;
      RECT  14.95 5.2 16.23 5.205 ;
      RECT  14.95 5.205 16.225 5.21 ;
      RECT  14.95 5.21 16.22 5.215 ;
      RECT  14.95 5.215 16.215 5.22 ;
      RECT  14.95 5.22 16.21 5.225 ;
      RECT  14.95 5.225 16.205 5.23 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.66 4.365 6.275 4.595 ;
      RECT  6.045 4.595 6.275 4.925 ;
      RECT  6.045 4.925 10.25 5.155 ;
      RECT  6.9 4.41 11.02 4.64 ;
      RECT  14.445 4.89 14.675 5.0 ;
      RECT  12.71 5.0 14.675 5.23 ;
      RECT  2.63 5.0 5.21 5.23 ;
      RECT  19.43 5.0 21.45 5.23 ;
  END
END MDN_FSDPHRBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDPHRBQ_4
#      Description : D-Flip Flop w/scan, pos-edge triggered, lo-async-clear, sync hold, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(iq&EN&!SE)|(!EN&(!SE&D))|(SE&SI),clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDPHRBQ_4
  CLASS CORE ;
  FOREIGN MDN_FSDPHRBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 31.36 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  29.51 0.37 29.85 0.6 ;
      RECT  29.54 0.6 29.82 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 2.1 8.515 2.38 ;
      RECT  8.285 2.38 8.515 2.69 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 11.9 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  24.12 1.565 27.4 1.795 ;
      RECT  26.765 1.795 26.995 3.245 ;
      RECT  24.12 3.245 27.4 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.22 2.125 18.62 2.355 ;
      RECT  17.22 2.355 17.5 2.915 ;
      RECT  18.34 2.355 18.62 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 2.94 2.355 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  30.125 4.9 30.355 5.46 ;
      RECT  30.125 5.46 31.53 5.74 ;
      RECT  27.885 4.87 28.115 5.46 ;
      RECT  27.885 5.46 28.56 5.74 ;
      RECT  25.645 4.87 25.875 5.46 ;
      RECT  25.645 5.46 26.32 5.74 ;
      RECT  23.405 4.87 23.635 5.46 ;
      RECT  22.96 5.46 23.635 5.74 ;
      RECT  18.925 4.985 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 5.08 16.915 5.46 ;
      RECT  16.24 5.46 17.36 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 31.36 5.74 ;
      LAYER VIA12 ;
      RECT  30.39 5.47 30.65 5.73 ;
      RECT  30.95 5.47 31.21 5.73 ;
      RECT  28.15 5.47 28.41 5.73 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  30.125 -0.14 31.53 0.14 ;
      RECT  30.125 0.14 30.355 0.7 ;
      RECT  25.645 -0.14 28.115 0.14 ;
      RECT  25.645 0.14 25.875 0.73 ;
      RECT  27.885 0.14 28.115 0.73 ;
      RECT  23.405 -0.14 24.08 0.14 ;
      RECT  23.405 0.14 23.635 0.52 ;
      RECT  17.36 -0.14 18.48 0.14 ;
      RECT  17.805 0.14 18.035 1.005 ;
      RECT  17.4 1.005 18.44 1.235 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 31.36 0.14 ;
      LAYER VIA12 ;
      RECT  30.39 -0.13 30.65 0.13 ;
      RECT  30.95 -0.13 31.21 0.13 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  27.03 -0.13 27.29 0.13 ;
      RECT  27.59 -0.13 27.85 0.13 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  18.07 -0.13 18.33 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  7.11 0.37 7.45 0.445 ;
      RECT  7.11 0.445 11.61 0.675 ;
      RECT  11.38 0.675 11.61 1.005 ;
      RECT  11.38 1.005 12.435 1.235 ;
      RECT  12.205 1.235 12.435 3.245 ;
      RECT  11.38 3.245 12.435 3.475 ;
      RECT  26.15 0.37 27.61 0.6 ;
      RECT  3.19 0.445 4.595 0.675 ;
      RECT  4.365 0.675 4.595 1.565 ;
      RECT  4.365 1.565 9.48 1.795 ;
      RECT  8.845 1.795 9.075 3.03 ;
      RECT  7.67 3.03 9.075 3.26 ;
      RECT  20.55 0.37 20.89 0.75 ;
      RECT  18.67 0.75 24.195 0.98 ;
      RECT  23.965 0.98 24.195 1.005 ;
      RECT  18.67 0.98 18.9 1.565 ;
      RECT  23.965 1.005 28.115 1.235 ;
      RECT  27.885 1.235 28.115 1.565 ;
      RECT  13.83 0.37 17.135 0.6 ;
      RECT  16.905 0.6 17.135 1.565 ;
      RECT  16.905 1.565 18.9 1.795 ;
      RECT  27.885 1.565 28.94 1.795 ;
      RECT  27.885 1.795 28.115 3.245 ;
      RECT  27.885 3.245 28.94 3.475 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 1.565 ;
      RECT  1.005 1.565 2.76 1.795 ;
      RECT  1.72 1.005 4.035 1.235 ;
      RECT  3.805 1.235 4.035 2.125 ;
      RECT  3.805 2.125 6.275 2.355 ;
      RECT  6.045 2.355 6.275 2.69 ;
      RECT  3.805 2.355 4.035 3.805 ;
      RECT  1.72 3.805 4.035 4.035 ;
      RECT  6.2 1.005 11.02 1.235 ;
      RECT  19.64 1.21 23.635 1.44 ;
      RECT  23.405 1.44 23.635 2.405 ;
      RECT  22.91 2.405 26.49 2.635 ;
      RECT  23.405 2.635 23.635 3.95 ;
      RECT  20.16 3.95 23.635 4.065 ;
      RECT  18.1 4.065 23.635 4.18 ;
      RECT  18.1 4.18 20.385 4.295 ;
      RECT  13.62 1.29 16.2 1.52 ;
      RECT  29.3 1.565 29.795 1.795 ;
      RECT  29.565 1.795 29.795 2.405 ;
      RECT  28.39 2.405 29.795 2.635 ;
      RECT  29.565 2.635 29.795 3.245 ;
      RECT  29.3 3.245 29.795 3.475 ;
      RECT  19.13 1.67 20.68 1.9 ;
      RECT  19.13 1.9 19.36 3.03 ;
      RECT  18.925 3.03 22.22 3.145 ;
      RECT  12.765 0.83 16.66 1.06 ;
      RECT  12.765 1.06 12.995 1.565 ;
      RECT  16.43 1.06 16.66 2.405 ;
      RECT  12.765 1.565 13.26 1.795 ;
      RECT  12.765 1.795 12.995 3.245 ;
      RECT  16.07 2.405 16.66 2.635 ;
      RECT  16.43 2.635 16.66 3.145 ;
      RECT  16.43 3.145 22.22 3.26 ;
      RECT  12.765 3.245 13.26 3.475 ;
      RECT  16.43 3.26 19.155 3.375 ;
      RECT  21.11 1.67 21.45 1.9 ;
      RECT  21.11 1.9 21.34 2.405 ;
      RECT  19.59 2.405 21.34 2.635 ;
      RECT  21.88 1.67 22.92 1.9 ;
      RECT  22.45 1.9 22.68 3.49 ;
      RECT  19.485 3.49 22.92 3.605 ;
      RECT  15.385 3.605 22.92 3.72 ;
      RECT  15.385 3.72 19.715 3.835 ;
      RECT  15.385 3.835 15.615 4.005 ;
      RECT  14.445 4.005 15.615 4.235 ;
      RECT  14.445 4.235 14.675 4.365 ;
      RECT  11.645 4.365 14.675 4.595 ;
      RECT  11.645 4.595 11.875 5.0 ;
      RECT  10.48 5.0 11.875 5.215 ;
      RECT  10.48 5.215 11.87 5.23 ;
      RECT  14.39 1.75 14.73 1.98 ;
      RECT  14.39 1.98 14.62 2.975 ;
      RECT  14.39 2.975 14.675 3.315 ;
      RECT  15.005 1.75 15.5 1.98 ;
      RECT  15.005 1.98 15.235 3.2 ;
      RECT  14.925 3.2 15.235 3.43 ;
      RECT  14.925 3.43 15.155 3.545 ;
      RECT  13.73 3.545 15.155 3.775 ;
      RECT  13.73 3.775 13.96 3.805 ;
      RECT  9.965 3.805 13.96 3.95 ;
      RECT  7.67 3.95 13.96 4.035 ;
      RECT  7.67 4.035 10.195 4.18 ;
      RECT  3.245 1.51 3.475 3.53 ;
      RECT  8.44 3.49 9.48 3.72 ;
      RECT  15.845 4.065 17.74 4.295 ;
      RECT  15.845 4.295 16.075 4.465 ;
      RECT  15.16 4.465 16.075 4.695 ;
      RECT  23.965 4.365 28.62 4.41 ;
      RECT  20.6 4.41 28.62 4.525 ;
      RECT  16.58 4.525 28.62 4.53 ;
      RECT  16.575 4.53 28.62 4.535 ;
      RECT  16.57 4.535 28.62 4.54 ;
      RECT  16.565 4.54 28.62 4.545 ;
      RECT  16.56 4.545 28.62 4.55 ;
      RECT  16.555 4.55 28.62 4.555 ;
      RECT  16.55 4.555 28.62 4.56 ;
      RECT  16.545 4.56 28.62 4.565 ;
      RECT  16.54 4.565 28.62 4.57 ;
      RECT  16.535 4.57 28.62 4.575 ;
      RECT  16.53 4.575 28.62 4.58 ;
      RECT  16.525 4.58 28.62 4.585 ;
      RECT  16.52 4.585 28.62 4.59 ;
      RECT  16.515 4.59 28.62 4.595 ;
      RECT  16.51 4.595 24.195 4.6 ;
      RECT  28.39 4.595 28.62 5.0 ;
      RECT  16.505 4.6 24.195 4.605 ;
      RECT  16.5 4.605 24.195 4.61 ;
      RECT  16.495 4.61 24.195 4.615 ;
      RECT  16.49 4.615 24.195 4.62 ;
      RECT  16.485 4.62 24.195 4.625 ;
      RECT  16.48 4.625 24.195 4.63 ;
      RECT  16.475 4.63 24.195 4.635 ;
      RECT  16.47 4.635 24.195 4.64 ;
      RECT  16.465 4.64 20.845 4.645 ;
      RECT  21.67 4.64 21.9 5.0 ;
      RECT  16.46 4.645 20.845 4.65 ;
      RECT  16.455 4.65 20.845 4.655 ;
      RECT  16.45 4.655 20.845 4.66 ;
      RECT  16.445 4.66 20.845 4.665 ;
      RECT  16.44 4.665 20.845 4.67 ;
      RECT  16.435 4.67 20.845 4.675 ;
      RECT  16.43 4.675 20.845 4.68 ;
      RECT  16.425 4.68 20.845 4.685 ;
      RECT  16.42 4.685 20.845 4.69 ;
      RECT  16.415 4.69 20.845 4.695 ;
      RECT  16.41 4.695 20.845 4.7 ;
      RECT  16.405 4.7 20.845 4.705 ;
      RECT  16.4 4.705 20.845 4.71 ;
      RECT  16.395 4.71 20.845 4.715 ;
      RECT  16.39 4.715 20.845 4.72 ;
      RECT  16.385 4.72 20.845 4.725 ;
      RECT  16.38 4.725 20.845 4.73 ;
      RECT  16.375 4.73 20.845 4.735 ;
      RECT  16.37 4.735 20.845 4.74 ;
      RECT  16.365 4.74 20.845 4.745 ;
      RECT  16.36 4.745 20.845 4.75 ;
      RECT  16.355 4.75 20.845 4.755 ;
      RECT  16.35 4.755 16.675 4.76 ;
      RECT  16.345 4.76 16.67 4.765 ;
      RECT  16.34 4.765 16.665 4.77 ;
      RECT  16.335 4.77 16.66 4.775 ;
      RECT  16.33 4.775 16.655 4.78 ;
      RECT  16.325 4.78 16.65 4.785 ;
      RECT  16.32 4.785 16.645 4.79 ;
      RECT  16.315 4.79 16.64 4.795 ;
      RECT  16.31 4.795 16.635 4.8 ;
      RECT  16.305 4.8 16.63 4.805 ;
      RECT  16.3 4.805 16.625 4.81 ;
      RECT  16.295 4.81 16.62 4.815 ;
      RECT  16.29 4.815 16.615 4.82 ;
      RECT  16.285 4.82 16.61 4.825 ;
      RECT  16.28 4.825 16.605 4.83 ;
      RECT  16.275 4.83 16.6 4.835 ;
      RECT  16.27 4.835 16.595 4.84 ;
      RECT  16.265 4.84 16.59 4.845 ;
      RECT  16.26 4.845 16.585 4.85 ;
      RECT  16.255 4.85 16.58 4.855 ;
      RECT  16.25 4.855 16.575 4.86 ;
      RECT  16.245 4.86 16.57 4.865 ;
      RECT  16.24 4.865 16.565 4.87 ;
      RECT  16.235 4.87 16.56 4.875 ;
      RECT  16.23 4.875 16.555 4.88 ;
      RECT  16.225 4.88 16.55 4.885 ;
      RECT  16.22 4.885 16.545 4.89 ;
      RECT  16.215 4.89 16.54 4.895 ;
      RECT  16.21 4.895 16.535 4.9 ;
      RECT  16.205 4.9 16.53 4.905 ;
      RECT  16.2 4.905 16.525 4.91 ;
      RECT  16.195 4.91 16.52 4.915 ;
      RECT  16.19 4.915 16.515 4.92 ;
      RECT  16.185 4.92 16.51 4.925 ;
      RECT  16.18 4.925 16.505 4.93 ;
      RECT  16.175 4.93 16.5 4.935 ;
      RECT  16.17 4.935 16.495 4.94 ;
      RECT  16.165 4.94 16.49 4.945 ;
      RECT  16.16 4.945 16.485 4.95 ;
      RECT  16.155 4.95 16.48 4.955 ;
      RECT  16.15 4.955 16.475 4.96 ;
      RECT  16.145 4.96 16.47 4.965 ;
      RECT  16.14 4.965 16.465 4.97 ;
      RECT  16.135 4.97 16.46 4.975 ;
      RECT  16.13 4.975 16.455 4.98 ;
      RECT  16.125 4.98 16.45 4.985 ;
      RECT  16.12 4.985 16.445 4.99 ;
      RECT  16.115 4.99 16.44 4.995 ;
      RECT  16.11 4.995 16.435 5.0 ;
      RECT  14.95 5.0 16.43 5.005 ;
      RECT  21.67 5.0 22.01 5.23 ;
      RECT  28.39 5.0 28.73 5.23 ;
      RECT  14.95 5.005 16.425 5.01 ;
      RECT  14.95 5.01 16.42 5.015 ;
      RECT  14.95 5.015 16.415 5.02 ;
      RECT  14.95 5.02 16.41 5.025 ;
      RECT  14.95 5.025 16.405 5.03 ;
      RECT  14.95 5.03 16.4 5.035 ;
      RECT  14.95 5.035 16.395 5.04 ;
      RECT  14.95 5.04 16.39 5.045 ;
      RECT  14.95 5.045 16.385 5.05 ;
      RECT  14.95 5.05 16.38 5.055 ;
      RECT  14.95 5.055 16.375 5.06 ;
      RECT  14.95 5.06 16.37 5.065 ;
      RECT  14.95 5.065 16.365 5.07 ;
      RECT  14.95 5.07 16.36 5.075 ;
      RECT  14.95 5.075 16.355 5.08 ;
      RECT  14.95 5.08 16.35 5.085 ;
      RECT  14.95 5.085 16.345 5.09 ;
      RECT  14.95 5.09 16.34 5.095 ;
      RECT  14.95 5.095 16.335 5.1 ;
      RECT  14.95 5.1 16.33 5.105 ;
      RECT  14.95 5.105 16.325 5.11 ;
      RECT  14.95 5.11 16.32 5.115 ;
      RECT  14.95 5.115 16.315 5.12 ;
      RECT  14.95 5.12 16.31 5.125 ;
      RECT  14.95 5.125 16.305 5.13 ;
      RECT  14.95 5.13 16.3 5.135 ;
      RECT  14.95 5.135 16.295 5.14 ;
      RECT  14.95 5.14 16.29 5.145 ;
      RECT  14.95 5.145 16.285 5.15 ;
      RECT  14.95 5.15 16.28 5.155 ;
      RECT  14.95 5.155 16.275 5.16 ;
      RECT  14.95 5.16 16.27 5.165 ;
      RECT  14.95 5.165 16.265 5.17 ;
      RECT  14.95 5.17 16.26 5.175 ;
      RECT  14.95 5.175 16.255 5.18 ;
      RECT  14.95 5.18 16.25 5.185 ;
      RECT  14.95 5.185 16.245 5.19 ;
      RECT  14.95 5.19 16.24 5.195 ;
      RECT  14.95 5.195 16.235 5.2 ;
      RECT  14.95 5.2 16.23 5.205 ;
      RECT  14.95 5.205 16.225 5.21 ;
      RECT  14.95 5.21 16.22 5.215 ;
      RECT  14.95 5.215 16.215 5.22 ;
      RECT  14.95 5.22 16.21 5.225 ;
      RECT  14.95 5.225 16.205 5.23 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.66 4.365 6.275 4.595 ;
      RECT  6.045 4.595 6.275 4.925 ;
      RECT  6.045 4.925 10.25 5.155 ;
      RECT  6.9 4.41 11.02 4.64 ;
      RECT  14.445 4.89 14.675 5.0 ;
      RECT  12.71 5.0 14.675 5.23 ;
      RECT  21.165 4.89 21.395 5.0 ;
      RECT  19.43 5.0 21.395 5.23 ;
      RECT  2.63 5.0 5.21 5.23 ;
  END
END MDN_FSDPHRBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDPQ_1
#      Description : D-Flip Flop w/scan, pos-edge triggered, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDPQ_1
  CLASS CORE ;
  FOREIGN MDN_FSDPQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.245 1.565 17.74 1.795 ;
      RECT  17.245 1.795 17.475 3.245 ;
      RECT  17.245 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 12.435 5.74 ;
      RECT  12.205 5.0 12.435 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.6 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.36 -0.14 4.035 0.14 ;
      RECT  3.805 0.14 4.035 0.89 ;
      RECT  3.805 0.89 4.3 1.12 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  6.1 0.6 6.33 0.83 ;
      RECT  6.1 0.83 9.635 1.005 ;
      RECT  6.1 1.005 12.435 1.06 ;
      RECT  9.405 1.06 12.435 1.235 ;
      RECT  12.205 1.235 12.435 1.75 ;
      RECT  12.205 1.75 13.96 1.98 ;
      RECT  12.205 1.98 12.435 3.16 ;
      RECT  11.38 3.16 12.435 3.39 ;
      RECT  12.205 3.39 12.435 3.62 ;
      RECT  12.205 3.62 14.115 3.805 ;
      RECT  12.205 3.805 15.5 3.85 ;
      RECT  13.885 3.85 15.5 4.035 ;
      RECT  7.11 0.37 9.69 0.6 ;
      RECT  14.39 0.37 16.41 0.6 ;
      RECT  17.19 0.37 17.53 0.6 ;
      RECT  17.19 0.6 17.42 0.83 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.82 0.6 13.05 0.83 ;
      RECT  12.82 0.83 17.42 1.06 ;
      RECT  16.125 1.06 16.355 1.565 ;
      RECT  15.86 1.565 16.355 1.795 ;
      RECT  16.125 1.795 16.355 3.245 ;
      RECT  15.86 3.245 16.355 3.475 ;
      RECT  4.745 1.005 5.715 1.01 ;
      RECT  4.74 1.01 5.715 1.015 ;
      RECT  4.735 1.015 5.715 1.02 ;
      RECT  4.73 1.02 5.715 1.025 ;
      RECT  4.725 1.025 5.715 1.03 ;
      RECT  4.72 1.03 5.715 1.035 ;
      RECT  4.715 1.035 5.715 1.04 ;
      RECT  4.71 1.04 5.715 1.045 ;
      RECT  4.705 1.045 5.715 1.05 ;
      RECT  4.7 1.05 5.715 1.055 ;
      RECT  4.695 1.055 5.715 1.06 ;
      RECT  4.69 1.06 5.715 1.065 ;
      RECT  4.685 1.065 5.715 1.07 ;
      RECT  4.68 1.07 5.715 1.075 ;
      RECT  4.675 1.075 5.715 1.08 ;
      RECT  4.67 1.08 5.715 1.085 ;
      RECT  4.665 1.085 5.715 1.09 ;
      RECT  4.66 1.09 5.715 1.095 ;
      RECT  4.655 1.095 5.715 1.1 ;
      RECT  4.65 1.1 5.715 1.105 ;
      RECT  4.645 1.105 5.715 1.11 ;
      RECT  4.64 1.11 5.715 1.115 ;
      RECT  4.635 1.115 5.715 1.12 ;
      RECT  4.63 1.12 5.715 1.125 ;
      RECT  4.625 1.125 5.715 1.13 ;
      RECT  4.62 1.13 5.715 1.135 ;
      RECT  4.615 1.135 5.715 1.14 ;
      RECT  4.61 1.14 5.715 1.145 ;
      RECT  4.605 1.145 5.715 1.15 ;
      RECT  4.6 1.15 5.715 1.155 ;
      RECT  4.595 1.155 5.715 1.16 ;
      RECT  4.59 1.16 5.715 1.165 ;
      RECT  4.585 1.165 5.715 1.17 ;
      RECT  4.58 1.17 5.715 1.175 ;
      RECT  4.575 1.175 5.715 1.18 ;
      RECT  4.57 1.18 5.715 1.185 ;
      RECT  4.565 1.185 5.715 1.19 ;
      RECT  4.56 1.19 5.715 1.195 ;
      RECT  4.555 1.195 5.715 1.2 ;
      RECT  4.55 1.2 5.715 1.205 ;
      RECT  4.545 1.205 5.715 1.21 ;
      RECT  4.54 1.21 5.715 1.215 ;
      RECT  4.535 1.215 5.715 1.22 ;
      RECT  4.53 1.22 5.715 1.225 ;
      RECT  4.525 1.225 5.715 1.23 ;
      RECT  4.52 1.23 5.715 1.235 ;
      RECT  4.515 1.235 4.84 1.24 ;
      RECT  5.485 1.235 5.715 1.75 ;
      RECT  4.51 1.24 4.835 1.245 ;
      RECT  4.505 1.245 4.83 1.25 ;
      RECT  4.5 1.25 4.825 1.255 ;
      RECT  4.495 1.255 4.82 1.26 ;
      RECT  4.49 1.26 4.815 1.265 ;
      RECT  4.485 1.265 4.81 1.27 ;
      RECT  4.48 1.27 4.805 1.275 ;
      RECT  4.475 1.275 4.8 1.28 ;
      RECT  4.47 1.28 4.795 1.285 ;
      RECT  4.465 1.285 4.79 1.29 ;
      RECT  4.46 1.29 4.785 1.295 ;
      RECT  4.455 1.295 4.78 1.3 ;
      RECT  4.45 1.3 4.775 1.305 ;
      RECT  4.445 1.305 4.77 1.31 ;
      RECT  4.44 1.31 4.765 1.315 ;
      RECT  4.435 1.315 4.76 1.32 ;
      RECT  4.43 1.32 4.755 1.325 ;
      RECT  4.425 1.325 4.75 1.33 ;
      RECT  4.42 1.33 4.745 1.335 ;
      RECT  4.415 1.335 4.74 1.34 ;
      RECT  4.41 1.34 4.735 1.345 ;
      RECT  4.405 1.345 4.73 1.35 ;
      RECT  4.4 1.35 4.725 1.355 ;
      RECT  4.395 1.355 4.72 1.36 ;
      RECT  4.39 1.36 4.715 1.365 ;
      RECT  4.385 1.365 4.71 1.37 ;
      RECT  4.38 1.37 4.705 1.375 ;
      RECT  4.375 1.375 4.7 1.38 ;
      RECT  4.37 1.38 4.695 1.385 ;
      RECT  4.365 1.385 4.69 1.39 ;
      RECT  4.36 1.39 4.685 1.395 ;
      RECT  4.355 1.395 4.68 1.4 ;
      RECT  4.35 1.4 4.675 1.405 ;
      RECT  4.345 1.405 4.67 1.41 ;
      RECT  4.34 1.41 4.665 1.415 ;
      RECT  4.335 1.415 4.66 1.42 ;
      RECT  4.33 1.42 4.655 1.425 ;
      RECT  4.325 1.425 4.65 1.43 ;
      RECT  4.32 1.43 4.645 1.435 ;
      RECT  4.315 1.435 4.64 1.44 ;
      RECT  4.31 1.44 4.635 1.445 ;
      RECT  4.305 1.445 4.63 1.45 ;
      RECT  4.3 1.45 4.625 1.455 ;
      RECT  4.295 1.455 4.62 1.46 ;
      RECT  4.29 1.46 4.615 1.465 ;
      RECT  4.285 1.465 4.61 1.47 ;
      RECT  4.28 1.47 4.605 1.475 ;
      RECT  4.275 1.475 4.6 1.48 ;
      RECT  4.27 1.48 4.595 1.485 ;
      RECT  4.265 1.485 4.59 1.49 ;
      RECT  4.26 1.49 4.585 1.495 ;
      RECT  4.255 1.495 4.58 1.5 ;
      RECT  4.25 1.5 4.575 1.505 ;
      RECT  4.245 1.505 4.57 1.51 ;
      RECT  4.24 1.51 4.565 1.515 ;
      RECT  4.235 1.515 4.56 1.52 ;
      RECT  4.23 1.52 4.555 1.525 ;
      RECT  4.225 1.525 4.55 1.53 ;
      RECT  4.22 1.53 4.545 1.535 ;
      RECT  4.215 1.535 4.54 1.54 ;
      RECT  4.21 1.54 4.535 1.545 ;
      RECT  4.205 1.545 4.53 1.55 ;
      RECT  4.2 1.55 4.525 1.555 ;
      RECT  4.195 1.555 4.52 1.56 ;
      RECT  4.19 1.56 4.515 1.565 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  3.245 1.565 4.51 1.57 ;
      RECT  3.245 1.57 4.505 1.575 ;
      RECT  3.245 1.575 4.5 1.58 ;
      RECT  3.245 1.58 4.495 1.585 ;
      RECT  3.245 1.585 4.49 1.59 ;
      RECT  3.245 1.59 4.485 1.595 ;
      RECT  3.245 1.595 4.48 1.6 ;
      RECT  3.245 1.6 4.475 1.605 ;
      RECT  3.245 1.605 4.47 1.61 ;
      RECT  3.245 1.61 4.465 1.615 ;
      RECT  3.245 1.615 4.46 1.62 ;
      RECT  3.245 1.62 4.455 1.625 ;
      RECT  3.245 1.625 4.45 1.63 ;
      RECT  3.245 1.63 4.445 1.635 ;
      RECT  3.245 1.635 4.44 1.64 ;
      RECT  3.245 1.64 4.435 1.645 ;
      RECT  3.245 1.645 4.43 1.65 ;
      RECT  3.245 1.65 4.425 1.655 ;
      RECT  3.245 1.655 4.42 1.66 ;
      RECT  3.245 1.66 4.415 1.665 ;
      RECT  3.245 1.665 4.41 1.67 ;
      RECT  3.245 1.67 4.405 1.675 ;
      RECT  3.245 1.675 4.4 1.68 ;
      RECT  3.245 1.68 4.395 1.685 ;
      RECT  3.245 1.685 4.39 1.69 ;
      RECT  3.245 1.69 4.385 1.695 ;
      RECT  3.245 1.695 4.38 1.7 ;
      RECT  3.245 1.7 4.375 1.705 ;
      RECT  3.245 1.705 4.37 1.71 ;
      RECT  3.245 1.71 4.365 1.715 ;
      RECT  3.245 1.715 4.36 1.72 ;
      RECT  3.245 1.72 4.355 1.725 ;
      RECT  3.245 1.725 4.35 1.73 ;
      RECT  3.245 1.73 4.345 1.735 ;
      RECT  3.245 1.735 4.34 1.74 ;
      RECT  3.245 1.74 4.335 1.745 ;
      RECT  3.245 1.745 4.33 1.75 ;
      RECT  3.245 1.75 4.325 1.755 ;
      RECT  5.485 1.75 7.24 1.98 ;
      RECT  3.245 1.755 4.32 1.76 ;
      RECT  3.245 1.76 4.315 1.765 ;
      RECT  3.245 1.765 4.31 1.77 ;
      RECT  3.245 1.77 4.305 1.775 ;
      RECT  3.245 1.775 4.3 1.78 ;
      RECT  3.245 1.78 4.295 1.785 ;
      RECT  3.245 1.785 4.29 1.79 ;
      RECT  3.245 1.79 4.285 1.795 ;
      RECT  6.2 1.29 8.78 1.52 ;
      RECT  12.92 1.29 15.5 1.52 ;
      RECT  9.965 1.565 11.02 1.795 ;
      RECT  9.965 1.795 10.195 2.405 ;
      RECT  9.35 2.405 10.195 2.635 ;
      RECT  9.965 2.635 10.195 3.755 ;
      RECT  9.965 3.755 11.875 3.985 ;
      RECT  11.645 3.985 11.875 4.08 ;
      RECT  11.645 4.08 13.555 4.31 ;
      RECT  13.325 4.31 13.555 4.365 ;
      RECT  13.325 4.365 14.675 4.595 ;
      RECT  14.445 4.595 14.675 5.0 ;
      RECT  14.445 5.0 15.29 5.23 ;
      RECT  7.67 1.75 8.01 1.98 ;
      RECT  7.725 1.98 7.955 3.53 ;
      RECT  8.285 1.75 9.48 1.98 ;
      RECT  8.285 1.98 8.515 3.245 ;
      RECT  8.285 3.245 9.37 3.475 ;
      RECT  9.14 3.475 9.37 4.215 ;
      RECT  9.14 4.215 11.315 4.445 ;
      RECT  11.085 4.445 11.315 4.54 ;
      RECT  11.085 4.54 12.995 4.77 ;
      RECT  12.765 4.77 12.995 5.0 ;
      RECT  12.765 5.0 14.17 5.23 ;
      RECT  14.39 1.75 14.73 1.98 ;
      RECT  14.445 1.98 14.675 3.315 ;
      RECT  4.715 1.695 4.945 2.405 ;
      RECT  3.75 2.405 4.945 2.635 ;
      RECT  4.715 2.635 4.945 3.53 ;
      RECT  12.92 3.03 13.96 3.26 ;
      RECT  6.2 3.245 7.24 3.475 ;
      RECT  1.72 3.805 2.76 4.035 ;
      RECT  3.19 3.805 8.78 4.035 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  9.405 4.675 10.755 4.905 ;
      RECT  9.405 4.905 9.635 4.925 ;
      RECT  10.525 4.905 10.755 5.0 ;
      RECT  7.67 4.925 9.635 5.155 ;
      RECT  10.525 5.0 11.93 5.23 ;
      RECT  1.51 5.0 5.21 5.23 ;
  END
END MDN_FSDPQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDPQ_2
#      Description : D-Flip Flop w/scan, pos-edge triggered, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDPQ_2
  CLASS CORE ;
  FOREIGN MDN_FSDPQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.4 1.565 18.44 1.795 ;
      RECT  17.805 1.795 18.035 3.245 ;
      RECT  17.4 3.245 18.44 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 12.435 5.74 ;
      RECT  12.205 5.0 12.435 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 20.33 0.14 ;
      RECT  16.685 0.14 16.915 0.6 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  3.805 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.805 0.14 4.035 0.89 ;
      RECT  3.805 0.89 4.3 1.12 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  18.07 -0.13 18.33 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.98 0.37 6.32 0.375 ;
      RECT  5.98 0.375 6.46 0.6 ;
      RECT  6.23 0.6 6.46 0.83 ;
      RECT  6.23 0.83 9.62 1.005 ;
      RECT  6.23 1.005 12.435 1.06 ;
      RECT  9.39 1.06 12.435 1.235 ;
      RECT  12.205 1.235 12.435 1.75 ;
      RECT  12.205 1.75 13.96 1.98 ;
      RECT  12.205 1.98 12.435 3.16 ;
      RECT  11.38 3.16 12.435 3.39 ;
      RECT  12.205 3.39 12.435 3.62 ;
      RECT  12.205 3.62 14.115 3.805 ;
      RECT  12.205 3.805 15.5 3.85 ;
      RECT  13.885 3.85 15.5 4.035 ;
      RECT  7.11 0.37 9.69 0.6 ;
      RECT  14.39 0.37 16.41 0.6 ;
      RECT  17.19 0.37 18.65 0.6 ;
      RECT  17.19 0.6 17.42 0.83 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.82 0.6 13.05 0.83 ;
      RECT  12.82 0.83 17.42 1.06 ;
      RECT  16.125 1.06 16.355 1.565 ;
      RECT  15.86 1.565 16.355 1.795 ;
      RECT  16.125 1.795 16.355 3.245 ;
      RECT  15.86 3.245 16.355 3.475 ;
      RECT  4.745 1.005 5.715 1.01 ;
      RECT  4.74 1.01 5.715 1.015 ;
      RECT  4.735 1.015 5.715 1.02 ;
      RECT  4.73 1.02 5.715 1.025 ;
      RECT  4.725 1.025 5.715 1.03 ;
      RECT  4.72 1.03 5.715 1.035 ;
      RECT  4.715 1.035 5.715 1.04 ;
      RECT  4.71 1.04 5.715 1.045 ;
      RECT  4.705 1.045 5.715 1.05 ;
      RECT  4.7 1.05 5.715 1.055 ;
      RECT  4.695 1.055 5.715 1.06 ;
      RECT  4.69 1.06 5.715 1.065 ;
      RECT  4.685 1.065 5.715 1.07 ;
      RECT  4.68 1.07 5.715 1.075 ;
      RECT  4.675 1.075 5.715 1.08 ;
      RECT  4.67 1.08 5.715 1.085 ;
      RECT  4.665 1.085 5.715 1.09 ;
      RECT  4.66 1.09 5.715 1.095 ;
      RECT  4.655 1.095 5.715 1.1 ;
      RECT  4.65 1.1 5.715 1.105 ;
      RECT  4.645 1.105 5.715 1.11 ;
      RECT  4.64 1.11 5.715 1.115 ;
      RECT  4.635 1.115 5.715 1.12 ;
      RECT  4.63 1.12 5.715 1.125 ;
      RECT  4.625 1.125 5.715 1.13 ;
      RECT  4.62 1.13 5.715 1.135 ;
      RECT  4.615 1.135 5.715 1.14 ;
      RECT  4.61 1.14 5.715 1.145 ;
      RECT  4.605 1.145 5.715 1.15 ;
      RECT  4.6 1.15 5.715 1.155 ;
      RECT  4.595 1.155 5.715 1.16 ;
      RECT  4.59 1.16 5.715 1.165 ;
      RECT  4.585 1.165 5.715 1.17 ;
      RECT  4.58 1.17 5.715 1.175 ;
      RECT  4.575 1.175 5.715 1.18 ;
      RECT  4.57 1.18 5.715 1.185 ;
      RECT  4.565 1.185 5.715 1.19 ;
      RECT  4.56 1.19 5.715 1.195 ;
      RECT  4.555 1.195 5.715 1.2 ;
      RECT  4.55 1.2 5.715 1.205 ;
      RECT  4.545 1.205 5.715 1.21 ;
      RECT  4.54 1.21 5.715 1.215 ;
      RECT  4.535 1.215 5.715 1.22 ;
      RECT  4.53 1.22 5.715 1.225 ;
      RECT  4.525 1.225 5.715 1.23 ;
      RECT  4.52 1.23 5.715 1.235 ;
      RECT  4.515 1.235 4.84 1.24 ;
      RECT  5.485 1.235 5.715 1.75 ;
      RECT  4.51 1.24 4.835 1.245 ;
      RECT  4.505 1.245 4.83 1.25 ;
      RECT  4.5 1.25 4.825 1.255 ;
      RECT  4.495 1.255 4.82 1.26 ;
      RECT  4.49 1.26 4.815 1.265 ;
      RECT  4.485 1.265 4.81 1.27 ;
      RECT  4.48 1.27 4.805 1.275 ;
      RECT  4.475 1.275 4.8 1.28 ;
      RECT  4.47 1.28 4.795 1.285 ;
      RECT  4.465 1.285 4.79 1.29 ;
      RECT  4.46 1.29 4.785 1.295 ;
      RECT  4.455 1.295 4.78 1.3 ;
      RECT  4.45 1.3 4.775 1.305 ;
      RECT  4.445 1.305 4.77 1.31 ;
      RECT  4.44 1.31 4.765 1.315 ;
      RECT  4.435 1.315 4.76 1.32 ;
      RECT  4.43 1.32 4.755 1.325 ;
      RECT  4.425 1.325 4.75 1.33 ;
      RECT  4.42 1.33 4.745 1.335 ;
      RECT  4.415 1.335 4.74 1.34 ;
      RECT  4.41 1.34 4.735 1.345 ;
      RECT  4.405 1.345 4.73 1.35 ;
      RECT  4.4 1.35 4.725 1.355 ;
      RECT  4.395 1.355 4.72 1.36 ;
      RECT  4.39 1.36 4.715 1.365 ;
      RECT  4.385 1.365 4.71 1.37 ;
      RECT  4.38 1.37 4.705 1.375 ;
      RECT  4.375 1.375 4.7 1.38 ;
      RECT  4.37 1.38 4.695 1.385 ;
      RECT  4.365 1.385 4.69 1.39 ;
      RECT  4.36 1.39 4.685 1.395 ;
      RECT  4.355 1.395 4.68 1.4 ;
      RECT  4.35 1.4 4.675 1.405 ;
      RECT  4.345 1.405 4.67 1.41 ;
      RECT  4.34 1.41 4.665 1.415 ;
      RECT  4.335 1.415 4.66 1.42 ;
      RECT  4.33 1.42 4.655 1.425 ;
      RECT  4.325 1.425 4.65 1.43 ;
      RECT  4.32 1.43 4.645 1.435 ;
      RECT  4.315 1.435 4.64 1.44 ;
      RECT  4.31 1.44 4.635 1.445 ;
      RECT  4.305 1.445 4.63 1.45 ;
      RECT  4.3 1.45 4.625 1.455 ;
      RECT  4.295 1.455 4.62 1.46 ;
      RECT  4.29 1.46 4.615 1.465 ;
      RECT  4.285 1.465 4.61 1.47 ;
      RECT  4.28 1.47 4.605 1.475 ;
      RECT  4.275 1.475 4.6 1.48 ;
      RECT  4.27 1.48 4.595 1.485 ;
      RECT  4.265 1.485 4.59 1.49 ;
      RECT  4.26 1.49 4.585 1.495 ;
      RECT  4.255 1.495 4.58 1.5 ;
      RECT  4.25 1.5 4.575 1.505 ;
      RECT  4.245 1.505 4.57 1.51 ;
      RECT  4.24 1.51 4.565 1.515 ;
      RECT  4.235 1.515 4.56 1.52 ;
      RECT  4.23 1.52 4.555 1.525 ;
      RECT  4.225 1.525 4.55 1.53 ;
      RECT  4.22 1.53 4.545 1.535 ;
      RECT  4.215 1.535 4.54 1.54 ;
      RECT  4.21 1.54 4.535 1.545 ;
      RECT  4.205 1.545 4.53 1.55 ;
      RECT  4.2 1.55 4.525 1.555 ;
      RECT  4.195 1.555 4.52 1.56 ;
      RECT  4.19 1.56 4.515 1.565 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  3.245 1.565 4.51 1.57 ;
      RECT  3.245 1.57 4.505 1.575 ;
      RECT  3.245 1.575 4.5 1.58 ;
      RECT  3.245 1.58 4.495 1.585 ;
      RECT  3.245 1.585 4.49 1.59 ;
      RECT  3.245 1.59 4.485 1.595 ;
      RECT  3.245 1.595 4.48 1.6 ;
      RECT  3.245 1.6 4.475 1.605 ;
      RECT  3.245 1.605 4.47 1.61 ;
      RECT  3.245 1.61 4.465 1.615 ;
      RECT  3.245 1.615 4.46 1.62 ;
      RECT  3.245 1.62 4.455 1.625 ;
      RECT  3.245 1.625 4.45 1.63 ;
      RECT  3.245 1.63 4.445 1.635 ;
      RECT  3.245 1.635 4.44 1.64 ;
      RECT  3.245 1.64 4.435 1.645 ;
      RECT  3.245 1.645 4.43 1.65 ;
      RECT  3.245 1.65 4.425 1.655 ;
      RECT  3.245 1.655 4.42 1.66 ;
      RECT  3.245 1.66 4.415 1.665 ;
      RECT  3.245 1.665 4.41 1.67 ;
      RECT  3.245 1.67 4.405 1.675 ;
      RECT  3.245 1.675 4.4 1.68 ;
      RECT  3.245 1.68 4.395 1.685 ;
      RECT  3.245 1.685 4.39 1.69 ;
      RECT  3.245 1.69 4.385 1.695 ;
      RECT  3.245 1.695 4.38 1.7 ;
      RECT  3.245 1.7 4.375 1.705 ;
      RECT  3.245 1.705 4.37 1.71 ;
      RECT  3.245 1.71 4.365 1.715 ;
      RECT  3.245 1.715 4.36 1.72 ;
      RECT  3.245 1.72 4.355 1.725 ;
      RECT  3.245 1.725 4.35 1.73 ;
      RECT  3.245 1.73 4.345 1.735 ;
      RECT  3.245 1.735 4.34 1.74 ;
      RECT  3.245 1.74 4.335 1.745 ;
      RECT  3.245 1.745 4.33 1.75 ;
      RECT  3.245 1.75 4.325 1.755 ;
      RECT  5.485 1.75 7.24 1.98 ;
      RECT  3.245 1.755 4.32 1.76 ;
      RECT  3.245 1.76 4.315 1.765 ;
      RECT  3.245 1.765 4.31 1.77 ;
      RECT  3.245 1.77 4.305 1.775 ;
      RECT  3.245 1.775 4.3 1.78 ;
      RECT  3.245 1.78 4.295 1.785 ;
      RECT  3.245 1.785 4.29 1.79 ;
      RECT  3.245 1.79 4.285 1.795 ;
      RECT  6.2 1.29 8.78 1.52 ;
      RECT  12.92 1.29 15.5 1.52 ;
      RECT  9.965 1.565 11.02 1.795 ;
      RECT  9.965 1.795 10.195 2.405 ;
      RECT  9.35 2.405 10.195 2.635 ;
      RECT  9.965 2.635 10.195 3.755 ;
      RECT  9.965 3.755 11.875 3.985 ;
      RECT  11.645 3.985 11.875 4.08 ;
      RECT  11.645 4.08 13.555 4.31 ;
      RECT  13.325 4.31 13.555 4.52 ;
      RECT  13.325 4.52 14.675 4.75 ;
      RECT  14.445 4.75 14.675 5.0 ;
      RECT  14.445 5.0 15.29 5.23 ;
      RECT  4.66 1.75 5.155 1.98 ;
      RECT  4.925 1.98 5.155 2.405 ;
      RECT  3.75 2.405 5.155 2.635 ;
      RECT  4.925 2.635 5.155 3.245 ;
      RECT  4.66 3.245 5.155 3.475 ;
      RECT  7.67 1.75 8.01 1.98 ;
      RECT  7.725 1.98 7.955 3.435 ;
      RECT  8.285 1.75 9.485 1.98 ;
      RECT  8.285 1.98 8.515 3.245 ;
      RECT  8.285 3.245 9.635 3.475 ;
      RECT  9.405 3.475 9.635 4.215 ;
      RECT  9.14 4.215 11.315 4.445 ;
      RECT  11.085 4.445 11.315 4.54 ;
      RECT  11.085 4.54 12.995 4.77 ;
      RECT  12.765 4.77 12.995 5.0 ;
      RECT  12.765 5.0 14.17 5.23 ;
      RECT  14.39 1.75 14.73 1.98 ;
      RECT  14.445 1.98 14.675 3.315 ;
      RECT  12.92 3.16 13.96 3.39 ;
      RECT  6.2 3.245 7.24 3.475 ;
      RECT  1.72 3.805 2.76 4.035 ;
      RECT  3.19 3.805 8.78 4.035 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  9.405 4.675 10.75 4.905 ;
      RECT  9.405 4.905 9.635 4.925 ;
      RECT  10.52 4.905 10.75 5.0 ;
      RECT  7.67 4.925 9.635 5.155 ;
      RECT  10.52 5.0 11.93 5.23 ;
      RECT  1.51 5.0 5.21 5.23 ;
  END
END MDN_FSDPQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDPSBQ_2
#      Description : D-Flip Flop w/scan, pos-edge triggered, lo-async-/set, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDPSBQ_2
  CLASS CORE ;
  FOREIGN MDN_FSDPSBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.54 0.6 1.82 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.64 1.565 20.68 1.795 ;
      RECT  20.045 1.795 20.275 3.245 ;
      RECT  19.64 3.245 20.68 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.98 2.125 17.5 2.355 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.87 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  14.39 5.135 14.73 5.46 ;
      RECT  14.0 5.46 17.36 5.74 ;
      RECT  16.63 5.135 16.97 5.46 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.19 5.135 3.53 5.46 ;
      RECT  2.8 5.46 3.92 5.74 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  15.12 -0.14 16.24 0.14 ;
      RECT  15.215 0.14 15.445 1.005 ;
      RECT  15.215 1.005 17.74 1.235 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.685 -0.14 3.36 0.14 ;
      RECT  2.685 0.14 2.915 1.005 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  7.11 0.37 7.45 0.445 ;
      RECT  7.11 0.445 9.635 0.675 ;
      RECT  9.405 0.675 9.635 1.005 ;
      RECT  9.405 1.005 11.205 1.235 ;
      RECT  10.975 1.235 11.205 2.375 ;
      RECT  10.975 2.375 13.05 2.605 ;
      RECT  10.975 2.605 11.205 3.245 ;
      RECT  10.68 3.245 11.205 3.475 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  19.43 0.37 20.89 0.6 ;
      RECT  19.43 0.6 19.66 1.005 ;
      RECT  16.07 0.37 16.41 0.445 ;
      RECT  16.07 0.445 18.595 0.675 ;
      RECT  18.365 0.675 18.595 1.005 ;
      RECT  18.1 1.005 19.66 1.235 ;
      RECT  18.925 1.235 19.155 4.365 ;
      RECT  18.1 4.365 19.155 4.595 ;
      RECT  11.645 0.445 14.985 0.675 ;
      RECT  11.645 0.675 11.875 0.95 ;
      RECT  14.755 0.675 14.985 1.565 ;
      RECT  11.435 0.95 11.875 1.29 ;
      RECT  14.755 1.565 16.2 1.795 ;
      RECT  3.245 1.005 8.78 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  1.72 1.565 3.475 1.795 ;
      RECT  12.92 1.005 14.115 1.235 ;
      RECT  13.885 1.235 14.115 1.985 ;
      RECT  13.885 1.985 14.455 1.99 ;
      RECT  13.885 1.99 14.46 1.995 ;
      RECT  13.885 1.995 14.465 2.0 ;
      RECT  13.885 2.0 14.47 2.005 ;
      RECT  13.885 2.005 14.475 2.01 ;
      RECT  13.885 2.01 14.48 2.015 ;
      RECT  13.885 2.015 14.485 2.02 ;
      RECT  13.885 2.02 14.49 2.025 ;
      RECT  13.885 2.025 14.495 2.03 ;
      RECT  13.885 2.03 14.5 2.035 ;
      RECT  13.885 2.035 14.505 2.04 ;
      RECT  13.885 2.04 14.51 2.045 ;
      RECT  13.885 2.045 14.515 2.05 ;
      RECT  13.885 2.05 14.52 2.055 ;
      RECT  13.885 2.055 14.525 2.06 ;
      RECT  13.885 2.06 14.53 2.065 ;
      RECT  13.885 2.065 14.535 2.07 ;
      RECT  13.885 2.07 14.54 2.075 ;
      RECT  13.885 2.075 14.545 2.08 ;
      RECT  13.885 2.08 14.55 2.085 ;
      RECT  13.885 2.085 14.555 2.09 ;
      RECT  13.885 2.09 14.56 2.095 ;
      RECT  13.885 2.095 14.565 2.1 ;
      RECT  13.885 2.1 14.57 2.105 ;
      RECT  13.885 2.105 14.575 2.11 ;
      RECT  13.885 2.11 14.58 2.115 ;
      RECT  13.885 2.115 14.585 2.12 ;
      RECT  13.885 2.12 14.59 2.125 ;
      RECT  13.885 2.125 14.595 2.13 ;
      RECT  13.885 2.13 14.6 2.135 ;
      RECT  13.885 2.135 14.605 2.14 ;
      RECT  13.885 2.14 14.61 2.145 ;
      RECT  13.885 2.145 14.615 2.15 ;
      RECT  13.885 2.15 14.62 2.155 ;
      RECT  13.885 2.155 14.625 2.16 ;
      RECT  13.885 2.16 14.63 2.165 ;
      RECT  13.885 2.165 14.635 2.17 ;
      RECT  13.885 2.17 14.64 2.175 ;
      RECT  13.885 2.175 14.645 2.18 ;
      RECT  13.885 2.18 14.65 2.185 ;
      RECT  13.885 2.185 14.655 2.19 ;
      RECT  13.885 2.19 14.66 2.195 ;
      RECT  13.885 2.195 14.665 2.2 ;
      RECT  13.885 2.2 14.67 2.205 ;
      RECT  13.885 2.205 14.675 2.215 ;
      RECT  14.35 2.215 14.675 2.22 ;
      RECT  14.355 2.22 14.675 2.225 ;
      RECT  14.36 2.225 14.675 2.23 ;
      RECT  14.365 2.23 14.675 2.235 ;
      RECT  14.37 2.235 14.675 2.24 ;
      RECT  14.375 2.24 14.675 2.245 ;
      RECT  14.38 2.245 14.675 2.25 ;
      RECT  14.385 2.25 14.675 2.255 ;
      RECT  14.39 2.255 14.675 2.26 ;
      RECT  14.395 2.26 14.675 2.265 ;
      RECT  14.4 2.265 14.675 2.27 ;
      RECT  14.405 2.27 14.675 2.275 ;
      RECT  14.41 2.275 14.675 2.28 ;
      RECT  14.415 2.28 14.675 2.285 ;
      RECT  14.42 2.285 14.675 2.29 ;
      RECT  14.425 2.29 14.675 2.295 ;
      RECT  14.43 2.295 14.675 2.3 ;
      RECT  14.435 2.3 14.675 2.305 ;
      RECT  14.44 2.305 14.675 2.31 ;
      RECT  14.445 2.31 14.675 3.755 ;
      RECT  13.125 3.755 15.5 3.985 ;
      RECT  13.125 3.985 13.355 4.005 ;
      RECT  12.205 4.005 13.355 4.235 ;
      RECT  12.205 4.235 12.435 4.365 ;
      RECT  9.405 4.365 12.435 4.595 ;
      RECT  9.405 4.595 9.635 4.925 ;
      RECT  5.99 4.925 9.635 5.155 ;
      RECT  5.99 5.155 6.33 5.23 ;
      RECT  4.365 1.565 5.0 1.795 ;
      RECT  4.365 1.795 4.595 3.755 ;
      RECT  1.005 3.755 5.0 3.985 ;
      RECT  1.005 3.985 1.235 4.365 ;
      RECT  0.49 4.365 1.235 4.595 ;
      RECT  0.49 4.595 0.72 5.0 ;
      RECT  0.38 5.0 0.72 5.23 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  8.28 1.565 10.745 1.795 ;
      RECT  8.28 1.795 8.51 2.35 ;
      RECT  10.515 1.795 10.745 2.69 ;
      RECT  8.28 2.35 8.515 2.69 ;
      RECT  8.28 2.69 8.51 3.245 ;
      RECT  8.28 3.245 9.48 3.475 ;
      RECT  12.15 1.565 13.555 1.795 ;
      RECT  13.325 1.795 13.555 2.835 ;
      RECT  12.205 2.835 13.555 3.065 ;
      RECT  12.205 3.065 12.435 3.315 ;
      RECT  13.83 2.445 14.17 2.675 ;
      RECT  13.94 2.675 14.17 3.295 ;
      RECT  12.665 3.295 14.17 3.525 ;
      RECT  12.665 3.525 12.895 3.545 ;
      RECT  11.645 3.545 12.895 3.775 ;
      RECT  11.645 3.775 11.875 3.805 ;
      RECT  7.725 1.51 7.955 3.805 ;
      RECT  7.725 3.805 11.875 4.035 ;
      RECT  0.18 3.245 2.76 3.475 ;
      RECT  5.485 3.805 7.24 4.035 ;
      RECT  5.485 4.035 5.715 4.365 ;
      RECT  4.925 4.365 5.715 4.595 ;
      RECT  4.925 4.595 5.155 4.675 ;
      RECT  2.685 4.675 5.155 4.905 ;
      RECT  2.685 4.905 2.915 4.925 ;
      RECT  0.95 4.925 2.915 5.155 ;
      RECT  1.72 4.215 4.3 4.445 ;
      RECT  13.585 4.215 17.74 4.445 ;
      RECT  13.585 4.445 13.815 4.465 ;
      RECT  12.92 4.465 13.815 4.695 ;
      RECT  6.2 4.365 8.78 4.595 ;
      RECT  14.19 4.675 17.475 4.68 ;
      RECT  14.185 4.68 17.475 4.685 ;
      RECT  14.18 4.685 17.475 4.69 ;
      RECT  14.175 4.69 17.475 4.695 ;
      RECT  14.17 4.695 17.475 4.7 ;
      RECT  14.165 4.7 17.475 4.705 ;
      RECT  14.16 4.705 17.475 4.71 ;
      RECT  14.155 4.71 17.475 4.715 ;
      RECT  14.15 4.715 17.475 4.72 ;
      RECT  14.145 4.72 17.475 4.725 ;
      RECT  14.14 4.725 17.475 4.73 ;
      RECT  14.135 4.73 17.475 4.735 ;
      RECT  14.13 4.735 17.475 4.74 ;
      RECT  14.125 4.74 17.475 4.745 ;
      RECT  14.12 4.745 17.475 4.75 ;
      RECT  14.115 4.75 17.475 4.755 ;
      RECT  14.11 4.755 17.475 4.76 ;
      RECT  14.105 4.76 17.475 4.765 ;
      RECT  14.1 4.765 17.475 4.77 ;
      RECT  14.095 4.77 17.475 4.775 ;
      RECT  14.09 4.775 17.475 4.78 ;
      RECT  14.085 4.78 17.475 4.785 ;
      RECT  14.08 4.785 17.475 4.79 ;
      RECT  14.075 4.79 17.475 4.795 ;
      RECT  14.07 4.795 17.475 4.8 ;
      RECT  14.065 4.8 17.475 4.805 ;
      RECT  14.06 4.805 17.475 4.81 ;
      RECT  14.055 4.81 17.475 4.815 ;
      RECT  14.05 4.815 17.475 4.82 ;
      RECT  14.045 4.82 17.475 4.825 ;
      RECT  14.04 4.825 17.475 4.83 ;
      RECT  14.035 4.83 17.475 4.835 ;
      RECT  14.03 4.835 17.475 4.84 ;
      RECT  14.025 4.84 17.475 4.845 ;
      RECT  14.02 4.845 17.475 4.85 ;
      RECT  14.015 4.85 17.475 4.855 ;
      RECT  14.01 4.855 17.475 4.86 ;
      RECT  14.005 4.86 17.475 4.865 ;
      RECT  14.0 4.865 17.475 4.87 ;
      RECT  13.995 4.87 17.475 4.875 ;
      RECT  13.99 4.875 17.475 4.88 ;
      RECT  13.985 4.88 17.475 4.885 ;
      RECT  13.98 4.885 17.475 4.89 ;
      RECT  13.975 4.89 17.475 4.895 ;
      RECT  13.97 4.895 17.475 4.9 ;
      RECT  13.965 4.9 17.475 4.905 ;
      RECT  13.96 4.905 14.285 4.91 ;
      RECT  17.245 4.905 17.475 5.0 ;
      RECT  13.955 4.91 14.28 4.915 ;
      RECT  13.95 4.915 14.275 4.92 ;
      RECT  13.945 4.92 14.27 4.925 ;
      RECT  12.15 4.925 14.265 4.93 ;
      RECT  12.15 4.93 14.26 4.935 ;
      RECT  12.15 4.935 14.255 4.94 ;
      RECT  12.15 4.94 14.25 4.945 ;
      RECT  12.15 4.945 14.245 4.95 ;
      RECT  12.15 4.95 14.24 4.955 ;
      RECT  12.15 4.955 14.235 4.96 ;
      RECT  12.15 4.96 14.23 4.965 ;
      RECT  12.15 4.965 14.225 4.97 ;
      RECT  12.15 4.97 14.22 4.975 ;
      RECT  12.15 4.975 14.215 4.98 ;
      RECT  12.15 4.98 14.21 4.985 ;
      RECT  12.15 4.985 14.205 4.99 ;
      RECT  12.15 4.99 14.2 4.995 ;
      RECT  12.15 4.995 14.195 5.0 ;
      RECT  12.15 5.0 14.19 5.005 ;
      RECT  17.245 5.0 18.65 5.23 ;
      RECT  12.15 5.005 14.185 5.01 ;
      RECT  12.15 5.01 14.18 5.015 ;
      RECT  12.15 5.015 14.175 5.02 ;
      RECT  12.15 5.02 14.17 5.025 ;
      RECT  12.15 5.025 14.165 5.03 ;
      RECT  12.15 5.03 14.16 5.035 ;
      RECT  12.15 5.035 14.155 5.04 ;
      RECT  12.15 5.04 14.15 5.045 ;
      RECT  12.15 5.045 14.145 5.05 ;
      RECT  12.15 5.05 14.14 5.055 ;
      RECT  12.15 5.055 14.135 5.06 ;
      RECT  12.15 5.06 14.13 5.065 ;
      RECT  12.15 5.065 14.125 5.07 ;
      RECT  12.15 5.07 14.12 5.075 ;
      RECT  12.15 5.075 14.115 5.08 ;
      RECT  12.15 5.08 14.11 5.085 ;
      RECT  12.15 5.085 14.105 5.09 ;
      RECT  12.15 5.09 14.1 5.095 ;
      RECT  12.15 5.095 14.095 5.1 ;
      RECT  12.15 5.1 14.09 5.105 ;
      RECT  12.15 5.105 14.085 5.11 ;
      RECT  12.15 5.11 14.08 5.115 ;
      RECT  12.15 5.115 14.075 5.12 ;
      RECT  12.15 5.12 14.07 5.125 ;
      RECT  12.15 5.125 14.065 5.13 ;
      RECT  12.15 5.13 14.06 5.135 ;
      RECT  12.15 5.135 14.055 5.14 ;
      RECT  12.15 5.14 14.05 5.145 ;
      RECT  12.15 5.145 14.045 5.15 ;
      RECT  12.15 5.15 14.04 5.155 ;
      RECT  10.47 5.0 11.92 5.23 ;
  END
END MDN_FSDPSBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_FSDPSBQ_4
#      Description : D-Flip Flop w/scan, pos-edge triggered, lo-async-/set, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDPSBQ_4
  CLASS CORE ;
  FOREIGN MDN_FSDPSBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 24.64 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.54 0.6 1.82 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.64 1.565 22.92 1.795 ;
      RECT  22.285 1.795 22.515 3.245 ;
      RECT  19.64 3.245 22.92 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.98 2.125 17.5 2.355 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.81 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  20.72 5.46 21.395 5.74 ;
      RECT  18.925 4.87 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  14.39 5.135 14.73 5.46 ;
      RECT  14.0 5.46 17.36 5.74 ;
      RECT  16.63 5.135 16.97 5.46 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.19 5.135 3.53 5.46 ;
      RECT  2.8 5.46 3.92 5.74 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 24.64 5.74 ;
      LAYER VIA12 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  24.23 5.47 24.49 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 24.81 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  15.12 -0.14 16.24 0.14 ;
      RECT  15.215 0.14 15.445 1.005 ;
      RECT  15.215 1.005 17.74 1.235 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.685 -0.14 3.36 0.14 ;
      RECT  2.685 0.14 2.915 1.005 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 24.64 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  22.55 -0.13 22.81 0.13 ;
      RECT  23.11 -0.13 23.37 0.13 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  7.11 0.37 7.45 0.445 ;
      RECT  7.11 0.445 9.635 0.675 ;
      RECT  9.405 0.675 9.635 1.005 ;
      RECT  9.405 1.005 11.205 1.235 ;
      RECT  10.975 1.235 11.205 2.375 ;
      RECT  10.975 2.375 13.05 2.605 ;
      RECT  10.975 2.605 11.205 3.245 ;
      RECT  10.68 3.245 11.205 3.475 ;
      RECT  16.07 0.37 16.41 0.445 ;
      RECT  16.07 0.445 18.595 0.675 ;
      RECT  18.365 0.675 18.595 1.005 ;
      RECT  18.1 1.005 19.155 1.235 ;
      RECT  18.925 1.235 19.155 2.405 ;
      RECT  18.925 2.405 21.835 2.635 ;
      RECT  18.925 2.635 19.155 4.365 ;
      RECT  18.1 4.365 19.155 4.595 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  21.67 0.37 23.13 0.6 ;
      RECT  11.645 0.445 14.97 0.675 ;
      RECT  11.645 0.675 11.875 0.95 ;
      RECT  14.74 0.675 14.97 1.565 ;
      RECT  11.435 0.95 11.875 1.29 ;
      RECT  14.74 1.565 16.2 1.795 ;
      RECT  3.245 1.005 8.78 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  1.72 1.565 3.475 1.795 ;
      RECT  12.92 1.005 14.115 1.235 ;
      RECT  13.885 1.235 14.115 1.985 ;
      RECT  13.885 1.985 14.425 1.99 ;
      RECT  13.885 1.99 14.43 1.995 ;
      RECT  13.885 1.995 14.435 2.0 ;
      RECT  13.885 2.0 14.44 2.005 ;
      RECT  13.885 2.005 14.445 2.01 ;
      RECT  13.885 2.01 14.45 2.015 ;
      RECT  13.885 2.015 14.455 2.02 ;
      RECT  13.885 2.02 14.46 2.025 ;
      RECT  13.885 2.025 14.465 2.03 ;
      RECT  13.885 2.03 14.47 2.035 ;
      RECT  13.885 2.035 14.475 2.04 ;
      RECT  13.885 2.04 14.48 2.045 ;
      RECT  13.885 2.045 14.485 2.05 ;
      RECT  13.885 2.05 14.49 2.055 ;
      RECT  13.885 2.055 14.495 2.06 ;
      RECT  13.885 2.06 14.5 2.065 ;
      RECT  13.885 2.065 14.505 2.07 ;
      RECT  13.885 2.07 14.51 2.075 ;
      RECT  13.885 2.075 14.515 2.08 ;
      RECT  13.885 2.08 14.52 2.085 ;
      RECT  13.885 2.085 14.525 2.09 ;
      RECT  13.885 2.09 14.53 2.095 ;
      RECT  13.885 2.095 14.535 2.1 ;
      RECT  13.885 2.1 14.54 2.105 ;
      RECT  13.885 2.105 14.545 2.11 ;
      RECT  13.885 2.11 14.55 2.115 ;
      RECT  13.885 2.115 14.555 2.12 ;
      RECT  13.885 2.12 14.56 2.125 ;
      RECT  13.885 2.125 14.565 2.13 ;
      RECT  13.885 2.13 14.57 2.135 ;
      RECT  13.885 2.135 14.575 2.14 ;
      RECT  13.885 2.14 14.58 2.145 ;
      RECT  13.885 2.145 14.585 2.15 ;
      RECT  13.885 2.15 14.59 2.155 ;
      RECT  13.885 2.155 14.595 2.16 ;
      RECT  13.885 2.16 14.6 2.165 ;
      RECT  13.885 2.165 14.605 2.17 ;
      RECT  13.885 2.17 14.61 2.175 ;
      RECT  13.885 2.175 14.615 2.18 ;
      RECT  13.885 2.18 14.62 2.185 ;
      RECT  13.885 2.185 14.625 2.19 ;
      RECT  13.885 2.19 14.63 2.195 ;
      RECT  13.885 2.195 14.635 2.2 ;
      RECT  13.885 2.2 14.64 2.205 ;
      RECT  13.885 2.205 14.645 2.21 ;
      RECT  13.885 2.21 14.65 2.215 ;
      RECT  14.32 2.215 14.655 2.22 ;
      RECT  14.325 2.22 14.66 2.225 ;
      RECT  14.33 2.225 14.665 2.23 ;
      RECT  14.335 2.23 14.67 2.235 ;
      RECT  14.34 2.235 14.675 2.24 ;
      RECT  14.345 2.24 14.675 2.245 ;
      RECT  14.35 2.245 14.675 2.25 ;
      RECT  14.355 2.25 14.675 2.255 ;
      RECT  14.36 2.255 14.675 2.26 ;
      RECT  14.365 2.26 14.675 2.265 ;
      RECT  14.37 2.265 14.675 2.27 ;
      RECT  14.375 2.27 14.675 2.275 ;
      RECT  14.38 2.275 14.675 2.28 ;
      RECT  14.385 2.28 14.675 2.285 ;
      RECT  14.39 2.285 14.675 2.29 ;
      RECT  14.395 2.29 14.675 2.295 ;
      RECT  14.4 2.295 14.675 2.3 ;
      RECT  14.405 2.3 14.675 2.305 ;
      RECT  14.41 2.305 14.675 2.31 ;
      RECT  14.415 2.31 14.675 2.315 ;
      RECT  14.42 2.315 14.675 2.32 ;
      RECT  14.425 2.32 14.675 2.325 ;
      RECT  14.43 2.325 14.675 2.33 ;
      RECT  14.435 2.33 14.675 2.335 ;
      RECT  14.44 2.335 14.675 2.34 ;
      RECT  14.445 2.34 14.675 3.755 ;
      RECT  13.125 3.755 15.5 3.985 ;
      RECT  13.125 3.985 13.355 4.02 ;
      RECT  12.205 4.02 13.355 4.25 ;
      RECT  12.205 4.25 12.435 4.365 ;
      RECT  9.405 4.365 12.435 4.595 ;
      RECT  9.405 4.595 9.635 4.925 ;
      RECT  5.99 4.925 9.635 5.155 ;
      RECT  5.99 5.155 6.33 5.23 ;
      RECT  4.365 1.565 5.0 1.795 ;
      RECT  4.365 1.795 4.595 3.755 ;
      RECT  1.005 3.755 5.0 3.985 ;
      RECT  1.005 3.985 1.235 4.365 ;
      RECT  0.49 4.365 1.235 4.595 ;
      RECT  0.49 4.595 0.72 5.0 ;
      RECT  0.38 5.0 0.72 5.23 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  8.285 1.565 10.745 1.795 ;
      RECT  10.515 1.795 10.745 2.69 ;
      RECT  8.285 1.795 8.515 3.245 ;
      RECT  8.285 3.245 9.48 3.475 ;
      RECT  12.15 1.565 13.555 1.795 ;
      RECT  13.325 1.795 13.555 2.835 ;
      RECT  12.205 2.835 13.555 3.065 ;
      RECT  12.205 3.065 12.435 3.315 ;
      RECT  13.83 2.445 14.17 2.675 ;
      RECT  13.94 2.675 14.17 3.295 ;
      RECT  12.665 3.295 14.17 3.525 ;
      RECT  12.665 3.525 12.895 3.545 ;
      RECT  11.645 3.545 12.895 3.775 ;
      RECT  11.645 3.775 11.875 3.805 ;
      RECT  7.725 1.51 7.955 3.805 ;
      RECT  7.725 3.805 11.875 4.035 ;
      RECT  0.18 3.245 2.76 3.475 ;
      RECT  5.485 3.805 7.24 4.035 ;
      RECT  5.485 4.035 5.715 4.365 ;
      RECT  4.925 4.365 5.715 4.595 ;
      RECT  4.925 4.595 5.155 4.675 ;
      RECT  2.685 4.675 5.155 4.905 ;
      RECT  2.685 4.905 2.915 4.925 ;
      RECT  0.95 4.925 2.915 5.155 ;
      RECT  1.72 4.215 4.3 4.445 ;
      RECT  13.585 4.215 17.74 4.445 ;
      RECT  13.585 4.445 13.815 4.48 ;
      RECT  12.92 4.48 13.815 4.71 ;
      RECT  6.2 4.365 8.78 4.595 ;
      RECT  14.19 4.675 17.475 4.68 ;
      RECT  14.185 4.68 17.475 4.685 ;
      RECT  14.18 4.685 17.475 4.69 ;
      RECT  14.175 4.69 17.475 4.695 ;
      RECT  14.17 4.695 17.475 4.7 ;
      RECT  14.165 4.7 17.475 4.705 ;
      RECT  14.16 4.705 17.475 4.71 ;
      RECT  14.155 4.71 17.475 4.715 ;
      RECT  14.15 4.715 17.475 4.72 ;
      RECT  14.145 4.72 17.475 4.725 ;
      RECT  14.14 4.725 17.475 4.73 ;
      RECT  14.135 4.73 17.475 4.735 ;
      RECT  14.13 4.735 17.475 4.74 ;
      RECT  14.125 4.74 17.475 4.745 ;
      RECT  14.12 4.745 17.475 4.75 ;
      RECT  14.115 4.75 17.475 4.755 ;
      RECT  14.11 4.755 17.475 4.76 ;
      RECT  14.105 4.76 17.475 4.765 ;
      RECT  14.1 4.765 17.475 4.77 ;
      RECT  14.095 4.77 17.475 4.775 ;
      RECT  14.09 4.775 17.475 4.78 ;
      RECT  14.085 4.78 17.475 4.785 ;
      RECT  14.08 4.785 17.475 4.79 ;
      RECT  14.075 4.79 17.475 4.795 ;
      RECT  14.07 4.795 17.475 4.8 ;
      RECT  14.065 4.8 17.475 4.805 ;
      RECT  14.06 4.805 17.475 4.81 ;
      RECT  14.055 4.81 17.475 4.815 ;
      RECT  14.05 4.815 17.475 4.82 ;
      RECT  14.045 4.82 17.475 4.825 ;
      RECT  14.04 4.825 17.475 4.83 ;
      RECT  14.035 4.83 17.475 4.835 ;
      RECT  14.03 4.835 17.475 4.84 ;
      RECT  14.025 4.84 17.475 4.845 ;
      RECT  14.02 4.845 17.475 4.85 ;
      RECT  14.015 4.85 17.475 4.855 ;
      RECT  14.01 4.855 17.475 4.86 ;
      RECT  14.005 4.86 17.475 4.865 ;
      RECT  14.0 4.865 17.475 4.87 ;
      RECT  13.995 4.87 17.475 4.875 ;
      RECT  13.99 4.875 17.475 4.88 ;
      RECT  13.985 4.88 17.475 4.885 ;
      RECT  13.98 4.885 17.475 4.89 ;
      RECT  13.975 4.89 17.475 4.895 ;
      RECT  13.97 4.895 17.475 4.9 ;
      RECT  13.965 4.9 17.475 4.905 ;
      RECT  13.96 4.905 14.285 4.91 ;
      RECT  17.245 4.905 17.475 5.0 ;
      RECT  13.955 4.91 14.28 4.915 ;
      RECT  13.95 4.915 14.275 4.92 ;
      RECT  13.945 4.92 14.27 4.925 ;
      RECT  13.94 4.925 14.265 4.93 ;
      RECT  13.935 4.93 14.26 4.935 ;
      RECT  13.93 4.935 14.255 4.94 ;
      RECT  12.15 4.94 14.25 4.945 ;
      RECT  12.15 4.945 14.245 4.95 ;
      RECT  12.15 4.95 14.24 4.955 ;
      RECT  12.15 4.955 14.235 4.96 ;
      RECT  12.15 4.96 14.23 4.965 ;
      RECT  12.15 4.965 14.225 4.97 ;
      RECT  12.15 4.97 14.22 4.975 ;
      RECT  12.15 4.975 14.215 4.98 ;
      RECT  12.15 4.98 14.21 4.985 ;
      RECT  12.15 4.985 14.205 4.99 ;
      RECT  12.15 4.99 14.2 4.995 ;
      RECT  12.15 4.995 14.195 5.0 ;
      RECT  12.15 5.0 14.19 5.005 ;
      RECT  17.245 5.0 18.65 5.23 ;
      RECT  12.15 5.005 14.185 5.01 ;
      RECT  12.15 5.01 14.18 5.015 ;
      RECT  12.15 5.015 14.175 5.02 ;
      RECT  12.15 5.02 14.17 5.025 ;
      RECT  12.15 5.025 14.165 5.03 ;
      RECT  12.15 5.03 14.16 5.035 ;
      RECT  12.15 5.035 14.155 5.04 ;
      RECT  12.15 5.04 14.15 5.045 ;
      RECT  12.15 5.045 14.145 5.05 ;
      RECT  12.15 5.05 14.14 5.055 ;
      RECT  12.15 5.055 14.135 5.06 ;
      RECT  12.15 5.06 14.13 5.065 ;
      RECT  12.15 5.065 14.125 5.07 ;
      RECT  12.15 5.07 14.12 5.075 ;
      RECT  12.15 5.075 14.115 5.08 ;
      RECT  12.15 5.08 14.11 5.085 ;
      RECT  12.15 5.085 14.105 5.09 ;
      RECT  12.15 5.09 14.1 5.095 ;
      RECT  12.15 5.095 14.095 5.1 ;
      RECT  12.15 5.1 14.09 5.105 ;
      RECT  12.15 5.105 14.085 5.11 ;
      RECT  12.15 5.11 14.08 5.115 ;
      RECT  12.15 5.115 14.075 5.12 ;
      RECT  12.15 5.12 14.07 5.125 ;
      RECT  12.15 5.125 14.065 5.13 ;
      RECT  12.15 5.13 14.06 5.135 ;
      RECT  12.15 5.135 14.055 5.14 ;
      RECT  12.15 5.14 14.05 5.145 ;
      RECT  12.15 5.145 14.045 5.15 ;
      RECT  12.15 5.15 14.04 5.155 ;
      RECT  12.15 5.155 14.035 5.16 ;
      RECT  12.15 5.16 14.03 5.165 ;
      RECT  12.15 5.165 14.025 5.17 ;
      RECT  10.47 5.0 11.92 5.23 ;
  END
END MDN_FSDPSBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_1
#      Description : Inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_1
  CLASS CORE ;
  FOREIGN MDN_INV_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.24 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.905 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 2.24 5.74 ;
      LAYER VIA12 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 2.24 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.565 1.235 1.795 ;
      RECT  1.005 1.795 1.235 3.805 ;
      RECT  0.18 3.805 1.235 4.035 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
END MDN_INV_1
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_12
#      Description : Inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_12
  CLASS CORE ;
  FOREIGN MDN_INV_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.66 ;
      RECT  9.38 2.66 10.78 2.685 ;
      RECT  10.5 2.125 10.78 2.66 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 10.78 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
      RECT  2.66 2.125 2.94 2.685 ;
      RECT  3.78 2.125 4.06 2.685 ;
      RECT  4.9 2.125 5.18 2.685 ;
      RECT  6.02 2.125 6.3 2.685 ;
      RECT  7.14 2.125 7.42 2.685 ;
      RECT  8.26 2.125 8.54 2.685 ;
    END
    ANTENNAGATEAREA 6.804 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.52 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.52 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.52 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.52 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.52 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.52 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.235 0.75 13.205 1.31 ;
      RECT  11.01 1.31 11.39 3.55 ;
      RECT  0.235 3.55 13.205 4.11 ;
    END
    ANTENNADIFFAREA 18.144 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  11.62 2.125 13.02 2.355 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
      RECT  10.47 5.0 11.93 5.23 ;
  END
END MDN_INV_12
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_16
#      Description : Inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_16
  CLASS CORE ;
  FOREIGN MDN_INV_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  16.125 4.365 17.475 4.595 ;
      RECT  16.125 4.595 16.355 5.0 ;
      RECT  17.245 4.595 17.475 5.0 ;
      RECT  13.885 4.365 15.235 4.595 ;
      RECT  13.885 4.595 14.115 5.0 ;
      RECT  15.005 4.595 15.235 5.0 ;
      RECT  11.645 4.365 12.995 4.595 ;
      RECT  11.645 4.595 11.875 5.0 ;
      RECT  12.765 4.595 12.995 5.0 ;
      RECT  9.405 4.365 10.755 4.595 ;
      RECT  9.405 4.595 9.635 5.0 ;
      RECT  10.525 4.595 10.755 5.0 ;
      RECT  7.165 4.365 8.515 4.595 ;
      RECT  7.165 4.595 7.395 5.0 ;
      RECT  8.285 4.595 8.515 5.0 ;
      RECT  4.925 4.365 6.275 4.595 ;
      RECT  4.925 4.595 5.155 5.0 ;
      RECT  6.045 4.595 6.275 5.0 ;
      RECT  2.685 4.365 4.035 4.595 ;
      RECT  2.685 4.595 2.915 5.0 ;
      RECT  3.805 4.595 4.035 5.0 ;
      RECT  0.445 4.365 1.795 4.595 ;
      RECT  0.445 4.595 0.675 5.0 ;
      RECT  1.565 4.595 1.795 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  1.51 5.0 2.97 5.23 ;
      RECT  3.75 5.0 5.21 5.23 ;
      RECT  5.99 5.0 7.45 5.23 ;
      RECT  8.23 5.0 9.69 5.23 ;
      RECT  10.47 5.0 11.93 5.23 ;
      RECT  12.71 5.0 14.17 5.23 ;
      RECT  14.95 5.0 16.41 5.23 ;
      RECT  17.19 5.0 17.53 5.23 ;
    END
    ANTENNAGATEAREA 9.072 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  11.76 -0.14 12.435 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  7.725 -0.14 10.195 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.565 17.74 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  13.325 1.795 13.555 3.245 ;
      RECT  0.18 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 24.192 ;
  END X
END MDN_INV_16
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_2
#      Description : Inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_2
  CLASS CORE ;
  FOREIGN MDN_INV_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.24 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 3.805 ;
      RECT  0.42 3.805 1.82 4.035 ;
      RECT  1.54 2.125 1.82 3.805 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.565 4.365 2.06 4.595 ;
      RECT  1.565 4.595 1.795 5.46 ;
      RECT  1.565 5.46 2.41 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 2.24 5.74 ;
      LAYER VIA12 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.565 -0.14 2.41 0.14 ;
      RECT  1.565 0.14 1.795 1.005 ;
      RECT  1.565 1.005 2.06 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 2.24 0.14 ;
      LAYER VIA12 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 1.51 1.235 3.53 ;
    END
    ANTENNADIFFAREA 2.566 ;
  END X
END MDN_INV_2
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_3
#      Description : Inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_3
  CLASS CORE ;
  FOREIGN MDN_INV_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.14 1.005 2.9 1.235 ;
      RECT  2.125 1.235 2.355 3.805 ;
      RECT  0.14 3.805 2.9 4.035 ;
    END
    ANTENNADIFFAREA 4.536 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 2.97 0.6 ;
  END
END MDN_INV_3
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_4
#      Description : Inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_4
  CLASS CORE ;
  FOREIGN MDN_INV_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.74 4.34 3.98 4.62 ;
      RECT  2.74 4.62 2.97 5.0 ;
      RECT  3.75 4.62 3.98 5.0 ;
      RECT  0.445 4.34 1.74 4.62 ;
      RECT  0.445 4.62 0.73 5.0 ;
      RECT  1.51 4.62 1.74 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  1.51 5.0 2.97 5.23 ;
      RECT  3.75 5.0 4.09 5.23 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 4.65 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 4.65 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.565 4.3 1.795 ;
      RECT  2.125 1.795 2.355 3.245 ;
      RECT  0.18 3.245 4.3 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
END MDN_INV_4
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_6
#      Description : Inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_6
  CLASS CORE ;
  FOREIGN MDN_INV_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 6.89 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 0.98 6.54 1.26 ;
      RECT  4.34 1.26 4.62 3.78 ;
      RECT  0.18 3.78 6.54 4.06 ;
    END
    ANTENNADIFFAREA 9.072 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.09 0.445 ;
      RECT  3.75 0.445 5.21 0.675 ;
      RECT  4.87 0.37 5.21 0.445 ;
      RECT  4.925 2.125 6.3 2.355 ;
      RECT  4.925 2.355 5.155 2.62 ;
      RECT  6.02 2.355 6.3 2.915 ;
  END
END MDN_INV_6
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_8
#      Description : Inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_8
  CLASS CORE ;
  FOREIGN MDN_INV_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.165 4.365 8.515 4.595 ;
      RECT  7.165 4.595 7.395 4.9 ;
      RECT  8.285 4.595 8.515 5.0 ;
      RECT  4.925 4.365 6.275 4.595 ;
      RECT  4.925 4.595 5.155 4.9 ;
      RECT  6.045 4.595 6.275 4.9 ;
      RECT  2.685 4.365 4.035 4.595 ;
      RECT  2.685 4.595 2.915 4.9 ;
      RECT  3.805 4.595 4.035 4.9 ;
      RECT  0.445 4.365 1.795 4.595 ;
      RECT  1.565 4.595 1.795 4.9 ;
      RECT  0.445 4.595 0.675 5.0 ;
      RECT  1.565 4.9 2.915 5.0 ;
      RECT  3.805 4.9 5.155 5.0 ;
      RECT  6.045 4.9 7.395 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  1.51 5.0 2.97 5.18 ;
      RECT  3.75 5.0 5.21 5.18 ;
      RECT  5.99 5.0 7.45 5.18 ;
      RECT  8.23 5.0 8.57 5.23 ;
      RECT  1.51 5.18 1.85 5.23 ;
      RECT  2.63 5.18 2.97 5.23 ;
      RECT  3.75 5.18 4.09 5.23 ;
      RECT  4.87 5.18 5.21 5.23 ;
      RECT  5.99 5.18 6.33 5.23 ;
      RECT  7.11 5.18 7.45 5.23 ;
    END
    ANTENNAGATEAREA 4.536 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 9.13 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 5.715 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.235 1.495 8.725 1.865 ;
      RECT  2.125 1.865 2.355 3.175 ;
      RECT  6.605 1.865 6.835 3.175 ;
      RECT  0.235 3.175 8.725 3.545 ;
    END
    ANTENNADIFFAREA 12.096 ;
  END X
END MDN_INV_8
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_AS_1
#      Description : Inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_AS_1
  CLASS CORE ;
  FOREIGN MDN_INV_AS_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 1.565 2.06 1.795 ;
      RECT  1.54 1.795 1.82 2.125 ;
      RECT  1.54 2.125 2.94 2.355 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNADIFFAREA 0.614 ;
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.905 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.905 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 4.65 0.14 ;
      RECT  3.245 0.14 3.475 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 3.245 ;
      RECT  1.72 3.245 3.475 3.475 ;
    END
    ANTENNADIFFAREA 2.41 ;
  END X
END MDN_INV_AS_1
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_AS_12
#      Description : Inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_AS_12
  CLASS CORE ;
  FOREIGN MDN_INV_AS_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 29.12 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.95 0.37 28.73 0.7 ;
      RECT  14.95 0.7 15.28 0.98 ;
      RECT  13.83 0.37 14.17 0.6 ;
      RECT  13.885 0.6 14.115 0.98 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.765 0.6 12.995 0.98 ;
      RECT  11.59 0.37 11.93 0.6 ;
      RECT  11.645 0.6 11.875 0.98 ;
      RECT  10.47 0.37 10.81 0.6 ;
      RECT  10.525 0.6 10.755 0.98 ;
      RECT  9.35 0.37 9.69 0.6 ;
      RECT  9.405 0.6 9.635 0.98 ;
      RECT  8.23 0.37 8.57 0.6 ;
      RECT  8.285 0.6 8.515 0.98 ;
      RECT  7.11 0.37 7.45 0.6 ;
      RECT  7.165 0.6 7.395 0.98 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  6.045 0.6 6.275 0.98 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.925 0.6 5.155 0.98 ;
      RECT  3.75 0.37 4.09 0.6 ;
      RECT  3.805 0.6 4.035 0.98 ;
      RECT  2.63 0.37 2.97 0.6 ;
      RECT  2.685 0.6 2.915 0.98 ;
      RECT  1.54 0.98 15.28 1.26 ;
      RECT  1.54 1.26 1.82 1.565 ;
      RECT  1.54 1.565 2.06 1.795 ;
      RECT  1.54 1.795 1.82 2.915 ;
    END
    ANTENNADIFFAREA 0.614 ;
    ANTENNAGATEAREA 14.175 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  28.445 4.365 28.94 4.595 ;
      RECT  28.445 4.595 28.675 5.46 ;
      RECT  28.445 5.46 29.29 5.74 ;
      RECT  27.06 4.365 27.555 4.595 ;
      RECT  27.325 4.595 27.555 5.46 ;
      RECT  26.88 5.46 27.555 5.74 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.2 5.46 25.875 5.74 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  22.96 5.46 23.635 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 21.395 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  -0.17 5.46 0.56 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 29.12 5.74 ;
      LAYER VIA12 ;
      RECT  28.71 5.47 28.97 5.73 ;
      RECT  27.03 5.47 27.29 5.73 ;
      RECT  25.35 5.47 25.61 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  20.31 5.47 20.57 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  28.56 -0.14 29.29 0.14 ;
      RECT  19.6 -0.14 20.72 0.14 ;
      RECT  12.205 -0.14 14.675 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  2.07 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 29.12 0.14 ;
      LAYER VIA12 ;
      RECT  28.71 -0.13 28.97 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  20.31 -0.13 20.57 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 15.725 2.215 ;
      RECT  2.42 2.215 3.17 2.38 ;
      RECT  15.075 2.215 15.725 2.825 ;
      RECT  15.075 2.825 28.21 3.385 ;
      RECT  2.11 3.385 28.21 3.475 ;
      RECT  2.11 3.475 15.725 4.035 ;
    END
    ANTENNADIFFAREA 28.596 ;
  END X
END MDN_INV_AS_12
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_AS_16
#      Description : Inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_AS_16
  CLASS CORE ;
  FOREIGN MDN_INV_AS_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 38.08 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.43 0.37 37.69 0.6 ;
      RECT  19.46 0.6 37.69 0.7 ;
      RECT  19.46 0.7 19.74 0.98 ;
      RECT  18.31 0.37 18.65 0.6 ;
      RECT  18.34 0.6 18.62 0.98 ;
      RECT  17.19 0.37 17.53 0.6 ;
      RECT  17.22 0.6 17.5 0.98 ;
      RECT  16.07 0.37 16.41 0.6 ;
      RECT  16.1 0.6 16.38 0.98 ;
      RECT  14.95 0.37 15.29 0.6 ;
      RECT  14.98 0.6 15.26 0.98 ;
      RECT  13.83 0.37 14.17 0.6 ;
      RECT  13.86 0.6 14.14 0.98 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.74 0.6 13.02 0.98 ;
      RECT  11.59 0.37 11.93 0.6 ;
      RECT  11.62 0.6 11.9 0.98 ;
      RECT  10.47 0.37 10.81 0.6 ;
      RECT  10.5 0.6 10.78 0.98 ;
      RECT  9.35 0.37 9.69 0.6 ;
      RECT  9.38 0.6 9.66 0.98 ;
      RECT  8.23 0.37 8.57 0.6 ;
      RECT  8.26 0.6 8.54 0.98 ;
      RECT  7.11 0.37 7.45 0.6 ;
      RECT  7.14 0.6 7.42 0.98 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  6.02 0.6 6.3 0.98 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.9 0.6 5.18 0.98 ;
      RECT  3.75 0.37 4.09 0.6 ;
      RECT  3.78 0.6 4.06 0.98 ;
      RECT  2.63 0.37 2.97 0.6 ;
      RECT  2.66 0.6 2.94 0.98 ;
      RECT  1.54 0.98 19.74 1.26 ;
      RECT  1.54 1.26 1.82 1.565 ;
      RECT  1.54 1.565 2.06 1.795 ;
      RECT  1.54 1.795 1.82 2.915 ;
    END
    ANTENNADIFFAREA 0.614 ;
    ANTENNAGATEAREA 18.711 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  37.405 4.365 37.9 4.595 ;
      RECT  37.405 4.595 37.635 5.46 ;
      RECT  37.405 5.46 38.25 5.74 ;
      RECT  36.02 4.365 36.515 4.595 ;
      RECT  36.285 4.595 36.515 5.46 ;
      RECT  35.84 5.46 36.515 5.74 ;
      RECT  34.605 4.9 34.835 5.46 ;
      RECT  34.16 5.46 34.835 5.74 ;
      RECT  32.365 4.9 32.595 5.46 ;
      RECT  31.92 5.46 32.595 5.74 ;
      RECT  30.125 4.9 30.355 5.46 ;
      RECT  29.68 5.46 30.355 5.74 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.645 5.46 28.115 5.74 ;
      RECT  27.885 4.9 28.115 5.46 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  22.96 5.46 23.635 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  20.72 5.46 21.395 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  -0.17 5.46 0.56 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 38.08 5.74 ;
      LAYER VIA12 ;
      RECT  37.67 5.47 37.93 5.73 ;
      RECT  35.99 5.47 36.25 5.73 ;
      RECT  34.31 5.47 34.57 5.73 ;
      RECT  32.07 5.47 32.33 5.73 ;
      RECT  29.83 5.47 30.09 5.73 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  27.03 5.47 27.29 5.73 ;
      RECT  27.59 5.47 27.85 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  37.52 -0.14 38.25 0.14 ;
      RECT  26.32 -0.14 27.44 0.14 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.695 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.695 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.695 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  12.205 0.14 12.435 0.695 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.695 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 38.08 0.14 ;
      LAYER VIA12 ;
      RECT  37.67 -0.13 37.93 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  27.03 -0.13 27.29 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.38 1.52 22.54 1.85 ;
      RECT  21.98 1.85 22.54 2.775 ;
      RECT  2.38 1.85 2.94 3.185 ;
      RECT  11.89 1.85 12.45 3.185 ;
      RECT  21.98 2.775 37.165 3.185 ;
      RECT  2.38 3.185 37.165 3.515 ;
    END
    ANTENNADIFFAREA 38.236 ;
  END X
END MDN_INV_AS_16
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_AS_2
#      Description : Inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_AS_2
  CLASS CORE ;
  FOREIGN MDN_INV_AS_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 1.565 2.06 1.795 ;
      RECT  1.54 1.795 1.82 2.915 ;
    END
    ANTENNADIFFAREA 0.614 ;
    ANTENNAGATEAREA 2.835 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 5.715 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  2.07 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 4.3 1.795 ;
      RECT  2.685 1.795 2.915 3.805 ;
      RECT  2.42 3.805 6.54 4.035 ;
    END
    ANTENNADIFFAREA 4.82 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.09 0.6 ;
      RECT  3.75 0.6 3.98 1.0 ;
      RECT  1.51 0.37 2.97 0.6 ;
      RECT  2.74 0.6 2.97 1.0 ;
      RECT  2.74 1.0 3.98 1.23 ;
      RECT  3.78 2.125 4.06 2.685 ;
      RECT  3.78 2.685 6.3 2.915 ;
      RECT  4.9 2.125 5.18 2.685 ;
      RECT  6.02 2.125 6.3 2.685 ;
  END
END MDN_INV_AS_2
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_AS_3
#      Description : Inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_AS_3
  CLASS CORE ;
  FOREIGN MDN_INV_AS_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 1.565 2.06 1.795 ;
      RECT  1.54 1.795 1.82 2.125 ;
      RECT  1.54 2.125 4.06 2.355 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNADIFFAREA 0.614 ;
    ANTENNAGATEAREA 3.969 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.905 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.905 7.955 5.46 ;
      RECT  3.245 4.905 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.695 ;
      RECT  5.485 0.14 5.715 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 5.0 1.795 ;
      RECT  4.365 1.795 4.595 3.805 ;
      RECT  2.42 3.805 8.78 4.035 ;
    END
    ANTENNADIFFAREA 7.23 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
  END
END MDN_INV_AS_3
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_AS_4
#      Description : Inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_AS_4
  CLASS CORE ;
  FOREIGN MDN_INV_AS_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.46 0.37 10.8 0.6 ;
      RECT  10.515 0.6 10.745 1.005 ;
      RECT  8.23 0.37 9.69 0.6 ;
      RECT  8.285 0.6 8.515 1.005 ;
      RECT  9.405 0.6 9.635 1.005 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  6.045 0.6 6.275 1.005 ;
      RECT  7.165 0.6 7.395 1.005 ;
      RECT  3.75 0.37 5.22 0.6 ;
      RECT  3.805 0.6 4.035 1.005 ;
      RECT  4.925 0.6 5.155 1.005 ;
      RECT  2.64 0.37 2.98 0.6 ;
      RECT  2.685 0.6 2.915 1.005 ;
      RECT  1.565 1.005 4.035 1.235 ;
      RECT  4.925 1.005 6.275 1.235 ;
      RECT  7.165 1.005 8.515 1.235 ;
      RECT  9.405 1.005 10.745 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.54 1.565 2.06 1.795 ;
      RECT  1.54 1.795 1.82 2.915 ;
    END
    ANTENNADIFFAREA 0.614 ;
    ANTENNAGATEAREA 5.103 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  -0.17 5.46 0.56 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 -0.14 11.37 0.14 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 6.835 1.795 ;
      RECT  6.605 1.795 6.835 3.805 ;
      RECT  2.42 3.805 11.02 4.035 ;
    END
    ANTENNADIFFAREA 9.64 ;
  END X
END MDN_INV_AS_4
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_AS_6
#      Description : Inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_AS_6
  CLASS CORE ;
  FOREIGN MDN_INV_AS_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.23 0.37 15.29 0.6 ;
      RECT  8.285 0.6 8.515 1.005 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  6.045 0.6 6.275 1.005 ;
      RECT  7.165 0.6 7.395 1.005 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  3.805 0.6 4.035 1.005 ;
      RECT  4.925 0.6 5.155 1.005 ;
      RECT  2.63 0.37 2.97 0.6 ;
      RECT  2.685 0.6 2.915 1.005 ;
      RECT  1.565 1.005 4.035 1.235 ;
      RECT  4.925 1.005 6.275 1.235 ;
      RECT  7.165 1.005 8.515 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.54 1.565 2.06 1.795 ;
      RECT  1.54 1.795 1.82 2.915 ;
    END
    ANTENNADIFFAREA 0.614 ;
    ANTENNAGATEAREA 7.371 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  -0.17 5.46 0.56 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  15.12 -0.14 15.85 0.14 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.395 1.515 9.125 1.845 ;
      RECT  8.795 1.845 9.125 3.755 ;
      RECT  2.395 3.755 15.525 4.085 ;
    END
    ANTENNADIFFAREA 14.46 ;
  END X
END MDN_INV_AS_6
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_AS_8
#      Description : Inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_AS_8
  CLASS CORE ;
  FOREIGN MDN_INV_AS_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.47 0.37 19.77 0.6 ;
      RECT  10.525 0.6 10.755 1.005 ;
      RECT  9.35 0.37 9.69 0.6 ;
      RECT  9.405 0.6 9.635 1.005 ;
      RECT  8.23 0.37 8.57 0.6 ;
      RECT  8.285 0.6 8.515 1.005 ;
      RECT  7.11 0.37 7.45 0.6 ;
      RECT  7.165 0.6 7.395 1.005 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  6.045 0.6 6.275 1.005 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.925 0.6 5.155 1.005 ;
      RECT  3.75 0.37 4.09 0.6 ;
      RECT  3.805 0.6 4.035 1.005 ;
      RECT  2.63 0.37 2.97 0.6 ;
      RECT  2.685 0.6 2.915 1.005 ;
      RECT  1.565 1.005 10.755 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.54 1.565 2.06 1.795 ;
      RECT  1.54 1.795 1.82 2.915 ;
    END
    ANTENNADIFFAREA 0.614 ;
    ANTENNAGATEAREA 9.639 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  -0.17 5.46 0.56 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  19.6 -0.14 20.33 0.14 ;
      RECT  7.725 -0.14 10.195 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.475 1.63 11.01 2.1 ;
      RECT  10.5 2.1 11.01 3.31 ;
      RECT  2.37 3.22 2.8 3.31 ;
      RECT  2.37 3.31 19.92 3.32 ;
      RECT  2.37 3.32 19.925 3.66 ;
      RECT  2.37 3.66 19.92 3.78 ;
    END
    ANTENNADIFFAREA 19.28 ;
  END X
END MDN_INV_AS_8
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_S_1
#      Description : Symmetric rise/fall time inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_S_1
  CLASS CORE ;
  FOREIGN MDN_INV_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.24 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.6 ;
      RECT  1.54 0.6 1.82 0.985 ;
      RECT  0.39 0.37 0.73 0.6 ;
      RECT  0.42 0.6 0.7 0.985 ;
      RECT  0.42 0.985 1.82 1.235 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  1.005 5.46 2.41 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 2.24 5.74 ;
      LAYER VIA12 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 2.24 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.565 0.675 1.795 ;
      RECT  0.445 1.795 0.675 3.805 ;
      RECT  0.18 3.805 2.06 4.035 ;
    END
    ANTENNADIFFAREA 2.41 ;
  END X
END MDN_INV_S_1
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_S_12
#      Description : Symmetric rise/fall time inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_S_12
  CLASS CORE ;
  FOREIGN MDN_INV_S_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 26.88 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  26.15 0.37 26.49 0.6 ;
      RECT  26.18 0.6 26.46 1.01 ;
      RECT  25.03 0.37 25.37 0.6 ;
      RECT  25.06 0.6 25.34 1.01 ;
      RECT  23.91 0.37 24.25 0.6 ;
      RECT  23.94 0.6 24.22 1.01 ;
      RECT  22.79 0.37 23.13 0.6 ;
      RECT  22.82 0.6 23.1 1.01 ;
      RECT  21.67 0.37 22.01 0.6 ;
      RECT  21.7 0.6 21.98 1.01 ;
      RECT  20.55 0.37 20.89 0.6 ;
      RECT  20.58 0.6 20.86 1.01 ;
      RECT  19.43 0.37 19.77 0.6 ;
      RECT  19.46 0.6 19.74 1.01 ;
      RECT  18.31 0.37 18.65 0.6 ;
      RECT  18.34 0.6 18.62 1.01 ;
      RECT  17.19 0.37 17.53 0.6 ;
      RECT  17.22 0.6 17.5 1.01 ;
      RECT  16.07 0.37 16.41 0.6 ;
      RECT  16.1 0.6 16.38 1.01 ;
      RECT  14.95 0.37 15.29 0.6 ;
      RECT  14.98 0.6 15.26 1.01 ;
      RECT  13.83 0.37 14.17 0.6 ;
      RECT  13.86 0.6 14.14 1.01 ;
      RECT  12.74 1.01 26.46 1.235 ;
      RECT  12.74 1.235 26.44 1.24 ;
      RECT  12.74 1.24 13.02 2.125 ;
      RECT  0.42 2.125 13.02 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 13.608 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 4.87 25.875 5.46 ;
      RECT  25.645 5.46 27.05 5.74 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.08 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  20.72 5.46 21.84 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.48 5.46 19.6 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 17.36 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 15.12 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.64 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.68 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 26.88 5.74 ;
      LAYER VIA12 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 -0.14 27.05 0.14 ;
      RECT  25.645 0.14 25.875 0.7 ;
      RECT  23.405 -0.14 24.08 0.14 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  21.165 -0.14 21.84 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.925 -0.14 19.6 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  13.27 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 26.88 0.14 ;
      LAYER VIA12 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.49 1.54 14.14 1.64 ;
      RECT  13.49 1.64 26.7 1.795 ;
      RECT  24.12 1.565 26.7 1.64 ;
      RECT  13.49 1.795 24.77 2.1 ;
      RECT  24.12 2.1 24.77 3.245 ;
      RECT  13.49 2.1 14.14 3.385 ;
      RECT  24.12 3.245 26.7 3.385 ;
      RECT  0.235 3.385 26.7 3.475 ;
      RECT  0.235 3.475 24.78 4.035 ;
    END
    ANTENNADIFFAREA 28.92 ;
  END X
END MDN_INV_S_12
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_S_16
#      Description : Symmetric rise/fall time inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_S_16
  CLASS CORE ;
  FOREIGN MDN_INV_S_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 35.84 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  35.11 0.37 35.45 0.6 ;
      RECT  35.14 0.6 35.42 1.005 ;
      RECT  33.99 0.37 34.33 0.6 ;
      RECT  34.02 0.6 34.3 1.005 ;
      RECT  32.87 0.37 33.21 0.6 ;
      RECT  32.9 0.6 33.18 1.005 ;
      RECT  31.75 0.37 32.09 0.6 ;
      RECT  31.78 0.6 32.06 1.005 ;
      RECT  30.63 0.37 30.97 0.6 ;
      RECT  30.66 0.6 30.94 1.005 ;
      RECT  29.51 0.37 29.85 0.6 ;
      RECT  29.54 0.6 29.82 1.005 ;
      RECT  28.39 0.37 28.73 0.6 ;
      RECT  28.42 0.6 28.7 1.005 ;
      RECT  27.27 0.37 27.61 0.6 ;
      RECT  27.3 0.6 27.58 1.005 ;
      RECT  26.15 0.37 26.49 0.6 ;
      RECT  26.18 0.6 26.46 1.005 ;
      RECT  25.03 0.37 25.37 0.6 ;
      RECT  25.06 0.6 25.34 1.005 ;
      RECT  23.91 0.37 24.25 0.6 ;
      RECT  23.94 0.6 24.22 1.005 ;
      RECT  22.79 0.37 23.13 0.6 ;
      RECT  22.82 0.6 23.1 1.005 ;
      RECT  21.67 0.37 22.01 0.6 ;
      RECT  21.7 0.6 21.98 1.005 ;
      RECT  20.55 0.37 20.89 0.6 ;
      RECT  20.58 0.6 20.86 1.005 ;
      RECT  19.43 0.37 19.77 0.6 ;
      RECT  19.46 0.6 19.74 1.005 ;
      RECT  18.31 0.37 18.65 0.6 ;
      RECT  18.34 0.6 18.62 1.005 ;
      RECT  17.22 1.005 35.42 1.235 ;
      RECT  17.22 1.235 17.5 2.125 ;
      RECT  0.42 2.125 17.5 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 18.144 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  34.605 4.87 34.835 5.46 ;
      RECT  34.605 5.46 36.01 5.74 ;
      RECT  32.365 4.9 32.595 5.46 ;
      RECT  32.365 5.46 33.04 5.74 ;
      RECT  30.125 4.9 30.355 5.46 ;
      RECT  30.125 5.46 30.8 5.74 ;
      RECT  27.885 4.9 28.115 5.46 ;
      RECT  27.885 5.46 28.56 5.74 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.645 5.46 26.32 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 23.635 5.74 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.63 5.135 16.97 5.46 ;
      RECT  16.24 5.46 17.36 5.74 ;
      RECT  14.39 5.135 14.73 5.46 ;
      RECT  14.0 5.46 15.12 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 12.88 5.74 ;
      RECT  12.15 5.135 12.49 5.46 ;
      RECT  7.67 5.135 8.01 5.46 ;
      RECT  7.28 5.46 8.4 5.74 ;
      RECT  5.43 5.135 5.77 5.46 ;
      RECT  5.04 5.46 6.16 5.74 ;
      RECT  3.19 5.135 3.53 5.46 ;
      RECT  2.8 5.46 3.92 5.74 ;
      RECT  0.95 5.135 1.29 5.46 ;
      RECT  -0.17 5.46 1.68 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 35.84 5.74 ;
      LAYER VIA12 ;
      RECT  34.87 5.47 35.13 5.73 ;
      RECT  35.43 5.47 35.69 5.73 ;
      RECT  32.63 5.47 32.89 5.73 ;
      RECT  30.39 5.47 30.65 5.73 ;
      RECT  28.15 5.47 28.41 5.73 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  22.55 5.47 22.81 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  34.605 -0.14 36.01 0.14 ;
      RECT  34.605 0.14 34.835 0.7 ;
      RECT  32.365 -0.14 33.04 0.14 ;
      RECT  32.365 0.14 32.595 0.7 ;
      RECT  30.125 -0.14 30.8 0.14 ;
      RECT  30.125 0.14 30.355 0.7 ;
      RECT  27.885 -0.14 28.56 0.14 ;
      RECT  27.885 0.14 28.115 0.7 ;
      RECT  25.645 -0.14 26.32 0.14 ;
      RECT  25.645 0.14 25.875 0.7 ;
      RECT  21.165 -0.14 23.635 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  23.405 0.14 23.635 0.7 ;
      RECT  18.925 -0.14 19.6 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  10.64 -0.14 11.76 0.14 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 35.84 0.14 ;
      LAYER VIA12 ;
      RECT  34.87 -0.13 35.13 0.13 ;
      RECT  35.43 -0.13 35.69 0.13 ;
      RECT  32.63 -0.13 32.89 0.13 ;
      RECT  30.39 -0.13 30.65 0.13 ;
      RECT  28.15 -0.13 28.41 0.13 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  22.55 -0.13 22.81 0.13 ;
      RECT  23.11 -0.13 23.37 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.11 1.54 35.66 1.87 ;
      RECT  18.11 1.87 18.85 2.935 ;
      RECT  24.54 1.87 25.01 3.195 ;
      RECT  30.99 1.87 31.46 3.195 ;
      RECT  17.78 2.935 18.85 3.195 ;
      RECT  17.78 3.195 35.66 3.5 ;
      RECT  0.235 3.5 35.66 3.525 ;
      RECT  0.235 3.525 18.29 4.115 ;
    END
    ANTENNADIFFAREA 38.56 ;
  END X
END MDN_INV_S_16
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_S_2
#      Description : Symmetric rise/fall time inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_S_2
  CLASS CORE ;
  FOREIGN MDN_INV_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 1.82 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 4.65 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  0.56 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      RECT  3.245 0.14 3.475 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.125 1.565 4.3 1.795 ;
      RECT  2.125 1.795 2.355 3.805 ;
      RECT  0.18 3.805 4.3 4.035 ;
    END
    ANTENNADIFFAREA 4.82 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.445 ;
      RECT  1.51 0.445 2.97 0.675 ;
      RECT  2.63 0.37 2.97 0.445 ;
      RECT  2.66 2.125 2.94 2.685 ;
      RECT  2.66 2.685 4.06 2.915 ;
      RECT  3.78 2.125 4.06 2.685 ;
  END
END MDN_INV_S_2
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_S_3
#      Description : Symmetric rise/fall time inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_S_3
  CLASS CORE ;
  FOREIGN MDN_INV_S_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 4.06 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
      RECT  2.66 2.125 2.94 2.685 ;
      RECT  3.78 2.125 4.06 2.685 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  0.56 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 4.595 1.235 ;
      RECT  4.365 1.235 4.595 3.805 ;
      RECT  0.18 3.805 6.54 4.035 ;
    END
    ANTENNADIFFAREA 7.23 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.09 0.445 ;
      RECT  3.75 0.445 5.21 0.675 ;
      RECT  4.87 0.37 5.21 0.445 ;
      RECT  4.9 2.125 5.18 2.685 ;
      RECT  4.9 2.685 6.3 2.915 ;
      RECT  6.02 2.125 6.3 2.685 ;
  END
END MDN_INV_S_3
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_S_4
#      Description : Symmetric rise/fall time inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_S_4
  CLASS CORE ;
  FOREIGN MDN_INV_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 6.3 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
      RECT  2.66 2.125 2.94 2.685 ;
      RECT  3.78 2.125 4.06 2.685 ;
      RECT  4.9 2.125 5.18 2.685 ;
      RECT  6.02 2.125 6.3 2.685 ;
    END
    ANTENNAGATEAREA 4.536 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  0.56 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 6.835 1.235 ;
      RECT  6.605 1.235 6.835 3.805 ;
      RECT  0.18 3.805 8.78 4.035 ;
    END
    ANTENNADIFFAREA 9.64 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.445 ;
      RECT  5.99 0.445 7.45 0.675 ;
      RECT  7.11 0.37 7.45 0.445 ;
      RECT  7.14 2.125 7.42 2.685 ;
      RECT  7.14 2.685 8.54 2.915 ;
      RECT  8.26 2.125 8.54 2.685 ;
  END
END MDN_INV_S_4
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_S_6
#      Description : Symmetric rise/fall time inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_S_6
  CLASS CORE ;
  FOREIGN MDN_INV_S_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 10.78 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
      RECT  2.66 2.125 2.94 2.685 ;
      RECT  3.78 2.125 4.06 2.685 ;
      RECT  4.9 2.125 5.18 2.685 ;
      RECT  6.02 2.125 6.3 2.685 ;
      RECT  7.14 2.125 7.42 2.685 ;
      RECT  8.26 2.125 8.54 2.685 ;
      RECT  9.38 2.125 9.66 2.685 ;
      RECT  10.5 2.125 10.78 2.685 ;
    END
    ANTENNAGATEAREA 6.804 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 13.61 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.54 13.26 1.82 ;
      RECT  11.06 1.82 11.34 3.78 ;
      RECT  0.18 3.78 13.26 4.06 ;
    END
    ANTENNADIFFAREA 14.46 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  10.47 0.37 10.81 0.445 ;
      RECT  10.47 0.445 11.93 0.675 ;
      RECT  11.59 0.37 11.93 0.445 ;
      RECT  11.7 0.675 11.93 1.005 ;
      RECT  11.7 1.005 12.94 1.235 ;
  END
END MDN_INV_S_6
#-----------------------------------------------------------------------
#      Cell        : MDN_INV_S_8
#      Description : Symmetric rise/fall time inverter
#      Equation    : X=!A
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_INV_S_8
  CLASS CORE ;
  FOREIGN MDN_INV_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 15.26 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
      RECT  2.66 2.125 2.94 2.685 ;
      RECT  3.78 2.125 4.06 2.685 ;
      RECT  4.9 2.125 5.18 2.685 ;
      RECT  6.02 2.125 6.3 2.685 ;
      RECT  7.14 2.125 7.42 2.685 ;
      RECT  8.26 2.125 8.54 2.685 ;
      RECT  9.38 2.125 9.66 2.685 ;
      RECT  10.5 2.125 10.78 2.685 ;
      RECT  11.62 2.125 11.9 2.685 ;
      RECT  12.74 2.125 13.02 2.685 ;
      RECT  13.86 2.125 14.14 2.685 ;
      RECT  14.98 2.125 15.26 2.685 ;
    END
    ANTENNAGATEAREA 9.072 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.705 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.705 ;
      RECT  8.79 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.705 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.14 0.935 15.865 1.305 ;
      RECT  15.495 1.305 15.865 1.495 ;
      RECT  15.495 1.495 17.74 1.865 ;
      RECT  16.615 1.865 16.985 3.735 ;
      RECT  0.18 3.735 17.74 4.105 ;
    END
    ANTENNADIFFAREA 19.28 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  17.19 0.37 17.53 0.6 ;
      RECT  17.19 0.6 17.42 1.005 ;
      RECT  14.95 0.37 16.41 0.6 ;
      RECT  16.18 0.6 16.41 1.005 ;
      RECT  16.18 1.005 17.42 1.235 ;
  END
END MDN_INV_S_8
#-----------------------------------------------------------------------
#      Cell        : MDN_LDNQ_4
#      Description : D-latch, neg-gate, q-only
#      Equation    : iq,iqn=latch(enable=!G,data_in=D):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDNQ_4
  CLASS CORE ;
  FOREIGN MDN_LDNQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.44 1.565 11.72 1.795 ;
      RECT  11.085 1.795 11.315 3.245 ;
      RECT  8.44 3.245 11.72 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.445 ;
      RECT  1.51 0.445 4.09 0.675 ;
      RECT  3.75 0.37 4.09 0.445 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.005 6.54 1.235 ;
      RECT  1.72 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 2.405 ;
      RECT  2.125 2.405 2.97 2.635 ;
      RECT  2.125 2.635 2.355 3.245 ;
      RECT  1.72 3.245 2.355 3.475 ;
      RECT  3.19 1.565 4.035 1.795 ;
      RECT  3.805 1.795 4.035 2.405 ;
      RECT  3.805 2.405 5.21 2.635 ;
      RECT  3.805 2.635 4.035 3.245 ;
      RECT  3.19 3.245 4.035 3.475 ;
      RECT  4.66 1.565 5.715 1.795 ;
      RECT  5.485 1.795 5.715 2.405 ;
      RECT  5.485 2.405 6.33 2.635 ;
      RECT  5.485 2.635 5.715 3.245 ;
      RECT  4.66 3.245 5.715 3.475 ;
      RECT  6.9 1.565 7.395 1.795 ;
      RECT  7.165 1.795 7.395 2.125 ;
      RECT  7.165 2.125 10.755 2.355 ;
      RECT  8.285 2.355 8.515 2.69 ;
      RECT  9.405 2.355 9.635 2.69 ;
      RECT  10.525 2.355 10.755 2.69 ;
      RECT  7.165 2.355 7.395 3.245 ;
      RECT  6.9 3.245 7.395 3.475 ;
      RECT  2.42 3.805 6.54 4.035 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  5.99 5.0 7.45 5.23 ;
      RECT  10.47 5.0 11.93 5.23 ;
  END
END MDN_LDNQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_LDNQ_1
#      Description : D-latch, neg-gate, q-only
#      Equation    : iq,iqn=latch(enable=!G,data_in=D):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDNQ_1
  CLASS CORE ;
  FOREIGN MDN_LDNQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.605 1.565 7.24 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  6.605 3.245 7.24 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.445 ;
      RECT  1.51 0.445 4.09 0.675 ;
      RECT  3.75 0.37 4.09 0.445 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.005 6.54 1.235 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
      RECT  4.66 1.565 5.715 1.795 ;
      RECT  5.485 1.795 5.715 2.405 ;
      RECT  5.485 2.405 6.33 2.635 ;
      RECT  5.485 2.635 5.715 3.245 ;
      RECT  4.66 3.245 5.715 3.475 ;
      RECT  3.245 1.51 3.475 2.685 ;
      RECT  3.245 2.685 5.155 2.915 ;
      RECT  4.925 2.35 5.155 2.685 ;
      RECT  3.245 2.915 3.475 3.53 ;
      RECT  2.42 3.805 6.54 4.035 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.98 4.365 6.275 4.595 ;
      RECT  4.98 4.595 5.21 5.0 ;
      RECT  6.045 4.595 6.275 5.0 ;
      RECT  4.87 5.0 5.21 5.23 ;
      RECT  6.045 5.0 7.45 5.23 ;
  END
END MDN_LDNQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_LDNQ_2
#      Description : D-latch, neg-gate, q-only
#      Equation    : iq,iqn=latch(enable=!G,data_in=D):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDNQ_2
  CLASS CORE ;
  FOREIGN MDN_LDNQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 8.78 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  6.9 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 9.13 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.445 ;
      RECT  1.51 0.445 4.09 0.675 ;
      RECT  3.75 0.37 4.09 0.445 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.005 6.54 1.235 ;
      RECT  1.72 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 2.405 ;
      RECT  2.125 2.405 2.97 2.635 ;
      RECT  2.125 2.635 2.355 3.245 ;
      RECT  1.72 3.245 2.355 3.475 ;
      RECT  4.66 1.565 5.715 1.795 ;
      RECT  5.485 1.795 5.715 2.405 ;
      RECT  5.485 2.405 6.33 2.635 ;
      RECT  5.485 2.635 5.715 3.245 ;
      RECT  4.66 3.245 5.715 3.475 ;
      RECT  3.245 1.505 3.475 2.685 ;
      RECT  3.245 2.685 5.155 2.915 ;
      RECT  4.925 2.35 5.155 2.685 ;
      RECT  3.245 2.915 3.475 3.53 ;
      RECT  2.42 3.805 6.54 4.035 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.98 4.365 8.46 4.595 ;
      RECT  4.98 4.595 5.21 5.0 ;
      RECT  7.22 4.595 7.45 5.0 ;
      RECT  8.23 4.595 8.46 5.0 ;
      RECT  4.87 5.0 5.21 5.23 ;
      RECT  7.11 5.0 7.45 5.23 ;
      RECT  8.23 5.0 8.57 5.23 ;
  END
END MDN_LDNQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_LDNRBQ_4
#      Description : D-latch, neg-gate, lo-async-clear, q-only
#      Equation    : iq,iqn=latch(enable=!G,data_in=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDNRBQ_4
  CLASS CORE ;
  FOREIGN MDN_LDNRBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 7.42 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.685 4.365 4.035 4.595 ;
      RECT  2.685 4.595 2.915 4.925 ;
      RECT  3.805 4.595 4.035 5.0 ;
      RECT  1.54 4.365 1.82 4.9 ;
      RECT  1.54 4.9 2.05 4.925 ;
      RECT  1.51 4.925 2.92 5.155 ;
      RECT  3.805 5.0 5.2 5.23 ;
      RECT  1.51 5.155 2.05 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.38 1.565 15.5 1.795 ;
      RECT  13.325 1.795 13.555 3.245 ;
      RECT  11.38 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.605 0.37 8.57 0.6 ;
      RECT  6.605 0.6 6.835 1.005 ;
      RECT  3.5 1.005 6.835 1.235 ;
      RECT  3.5 1.235 3.73 2.125 ;
      RECT  2.685 2.125 3.73 2.355 ;
      RECT  2.685 2.355 2.915 3.0 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.705 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  8.4 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  8.845 0.14 9.075 1.005 ;
      RECT  8.44 1.005 9.075 1.235 ;
      RECT  1.68 -0.14 2.8 0.14 ;
      RECT  2.125 0.14 2.355 1.005 ;
      RECT  2.125 1.005 2.76 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.445 ;
      RECT  3.04 0.445 6.33 0.675 ;
      RECT  3.04 0.675 3.27 1.565 ;
      RECT  1.565 1.565 3.27 1.795 ;
      RECT  1.565 1.795 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  12.71 0.37 14.17 0.6 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  9.14 1.565 9.635 1.795 ;
      RECT  9.405 1.795 9.635 3.805 ;
      RECT  9.14 3.805 9.635 3.81 ;
      RECT  6.045 3.245 7.955 3.475 ;
      RECT  6.045 3.475 6.275 3.49 ;
      RECT  7.725 3.475 7.955 3.81 ;
      RECT  4.03 2.355 4.26 2.685 ;
      RECT  4.03 2.685 5.155 2.915 ;
      RECT  4.925 2.915 5.155 3.49 ;
      RECT  4.925 3.49 6.275 3.72 ;
      RECT  7.725 3.81 9.635 4.04 ;
      RECT  9.405 4.04 9.635 4.365 ;
      RECT  9.405 4.365 10.755 4.595 ;
      RECT  10.525 4.595 10.755 5.0 ;
      RECT  10.47 5.0 10.81 5.23 ;
      RECT  10.735 1.51 10.965 2.125 ;
      RECT  10.735 2.125 12.995 2.355 ;
      RECT  11.645 2.355 11.875 2.69 ;
      RECT  12.765 2.355 12.995 2.69 ;
      RECT  10.735 2.355 10.965 3.53 ;
      RECT  13.885 2.125 15.235 2.355 ;
      RECT  13.885 2.355 14.115 2.69 ;
      RECT  15.005 2.355 15.235 2.69 ;
      RECT  5.485 1.51 5.715 3.03 ;
      RECT  5.43 3.03 5.77 3.26 ;
      RECT  3.96 3.245 4.595 3.475 ;
      RECT  4.365 3.475 4.595 3.95 ;
      RECT  4.365 3.95 6.54 4.18 ;
      RECT  6.805 3.805 7.24 4.035 ;
      RECT  6.805 4.035 7.035 4.41 ;
      RECT  4.66 4.41 7.035 4.64 ;
      RECT  7.265 4.365 9.075 4.595 ;
      RECT  7.265 4.595 7.495 4.985 ;
      RECT  8.845 4.595 9.075 5.0 ;
      RECT  5.43 4.985 7.495 5.215 ;
      RECT  8.845 5.0 9.69 5.23 ;
  END
END MDN_LDNRBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_LDNRBQ_1
#      Description : D-latch, neg-gate, lo-async-clear, q-only
#      Equation    : iq,iqn=latch(enable=!G,data_in=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDNRBQ_1
  CLASS CORE ;
  FOREIGN MDN_LDNRBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 7.42 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.685 4.365 4.035 4.595 ;
      RECT  2.685 4.595 2.915 4.925 ;
      RECT  3.805 4.595 4.035 4.925 ;
      RECT  1.54 4.365 1.82 4.9 ;
      RECT  1.54 4.9 2.05 4.925 ;
      RECT  1.51 4.925 2.915 5.155 ;
      RECT  3.805 4.925 5.2 5.155 ;
      RECT  1.51 5.155 2.05 5.23 ;
      RECT  4.86 5.155 5.2 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.525 1.565 11.02 1.795 ;
      RECT  10.525 1.795 10.755 3.245 ;
      RECT  10.525 3.245 11.02 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.165 0.37 8.57 0.6 ;
      RECT  7.165 0.6 7.395 1.005 ;
      RECT  3.5 1.005 7.395 1.235 ;
      RECT  3.5 1.235 3.73 2.125 ;
      RECT  2.685 2.125 3.73 2.355 ;
      RECT  2.685 2.355 2.915 3.0 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  8.4 -0.14 9.52 0.14 ;
      RECT  8.845 0.14 9.075 1.005 ;
      RECT  8.44 1.005 9.075 1.235 ;
      RECT  1.68 -0.14 2.8 0.14 ;
      RECT  2.125 0.14 2.355 1.005 ;
      RECT  2.125 1.005 2.76 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.445 ;
      RECT  3.04 0.445 6.33 0.675 ;
      RECT  3.04 0.675 3.27 1.565 ;
      RECT  1.565 1.565 3.27 1.795 ;
      RECT  1.565 1.795 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  9.14 1.565 9.635 1.795 ;
      RECT  9.405 1.795 9.635 3.805 ;
      RECT  6.045 3.245 7.955 3.475 ;
      RECT  6.045 3.475 6.275 3.49 ;
      RECT  7.725 3.475 7.955 3.805 ;
      RECT  4.03 2.345 4.26 2.685 ;
      RECT  4.03 2.685 5.155 2.915 ;
      RECT  4.925 2.915 5.155 3.49 ;
      RECT  4.925 3.49 6.275 3.72 ;
      RECT  7.725 3.805 9.635 4.035 ;
      RECT  5.485 1.51 5.715 3.03 ;
      RECT  5.43 3.03 5.77 3.26 ;
      RECT  3.955 3.805 4.595 3.95 ;
      RECT  3.955 3.95 6.54 4.035 ;
      RECT  4.365 4.035 6.54 4.18 ;
      RECT  6.77 3.805 7.24 4.035 ;
      RECT  6.77 4.035 7.0 4.465 ;
      RECT  4.66 4.465 7.0 4.695 ;
      RECT  7.265 4.365 10.7 4.595 ;
      RECT  7.265 4.595 7.495 4.925 ;
      RECT  9.46 4.595 9.69 5.0 ;
      RECT  10.47 4.595 10.7 5.0 ;
      RECT  5.43 4.925 7.495 5.155 ;
      RECT  9.35 5.0 9.69 5.23 ;
      RECT  10.47 5.0 10.81 5.23 ;
  END
END MDN_LDNRBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_LDNRBQ_2
#      Description : D-latch, neg-gate, lo-async-clear, q-only
#      Equation    : iq,iqn=latch(enable=!G,data_in=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDNRBQ_2
  CLASS CORE ;
  FOREIGN MDN_LDNRBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.925 2.125 6.305 2.355 ;
      RECT  4.925 2.355 5.155 2.69 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.14 1.565 11.02 1.795 ;
      RECT  9.965 1.795 10.195 3.245 ;
      RECT  9.14 3.245 11.02 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  5.79 0.37 6.33 0.445 ;
      RECT  1.005 0.445 6.33 0.675 ;
      RECT  1.005 0.675 1.235 1.565 ;
      RECT  0.42 1.565 1.235 1.795 ;
      RECT  0.42 1.795 0.7 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.43 5.135 5.77 5.46 ;
      RECT  5.04 5.46 6.16 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  6.55 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  6.605 0.14 6.835 1.005 ;
      RECT  6.2 1.005 6.835 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 10.81 0.6 ;
      RECT  10.47 0.6 10.7 1.005 ;
      RECT  8.23 0.37 9.71 0.6 ;
      RECT  8.23 0.6 8.46 1.005 ;
      RECT  9.48 0.6 9.71 1.005 ;
      RECT  7.725 1.005 8.46 1.235 ;
      RECT  9.48 1.005 10.7 1.235 ;
      RECT  7.725 1.235 7.955 3.705 ;
      RECT  3.245 1.54 3.475 3.03 ;
      RECT  3.24 3.03 5.715 3.26 ;
      RECT  5.485 3.26 5.715 3.705 ;
      RECT  5.485 3.705 7.955 3.935 ;
      RECT  6.2 3.7 6.54 3.705 ;
      RECT  1.715 1.005 2.76 1.235 ;
      RECT  3.96 1.005 5.0 1.235 ;
      RECT  3.805 1.565 7.4 1.795 ;
      RECT  3.805 1.795 4.035 2.72 ;
      RECT  7.165 1.795 7.395 3.245 ;
      RECT  6.9 3.245 7.395 3.475 ;
      RECT  8.285 1.565 8.78 1.795 ;
      RECT  8.285 1.795 8.515 4.215 ;
      RECT  4.51 4.215 8.78 4.445 ;
      RECT  4.51 4.445 4.74 4.54 ;
      RECT  1.565 4.54 4.74 4.77 ;
      RECT  1.565 4.77 1.795 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  2.42 3.51 5.0 3.74 ;
      RECT  4.015 3.97 4.245 4.08 ;
      RECT  1.72 4.08 4.245 4.31 ;
      RECT  4.97 4.675 6.275 4.905 ;
      RECT  4.97 4.905 5.2 5.0 ;
      RECT  6.045 4.905 6.275 5.0 ;
      RECT  2.63 5.0 5.2 5.23 ;
      RECT  6.045 5.0 7.45 5.23 ;
  END
END MDN_LDNRBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_LDNRBSBQ_1
#      Description : D-latch, neg-gate, lo-async-clear, lo-async-set, q-only
#      Equation    : iq,iqn=latch(enable=!G,data_in=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDNRBSBQ_1
  CLASS CORE ;
  FOREIGN MDN_LDNRBSBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.39 5.18 3.475 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 3.245 ;
      RECT  15.005 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.74 4.365 13.02 5.0 ;
      RECT  12.71 5.0 13.05 5.23 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.39 10.78 3.475 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.14 4.365 9.635 4.595 ;
      RECT  9.405 4.595 9.635 5.46 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 9.635 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.58 ;
      RECT  10.08 -0.14 10.755 0.14 ;
      RECT  10.525 0.14 10.755 0.89 ;
      RECT  10.525 0.89 11.02 1.12 ;
      RECT  5.485 -0.14 6.72 0.14 ;
      RECT  5.485 0.14 5.715 1.005 ;
      RECT  5.485 1.005 7.24 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 0.81 ;
      RECT  11.645 0.81 12.94 1.04 ;
      RECT  11.645 1.04 11.875 1.29 ;
      RECT  11.18 1.29 11.875 1.295 ;
      RECT  11.175 1.295 11.875 1.3 ;
      RECT  11.17 1.3 11.875 1.305 ;
      RECT  11.165 1.305 11.875 1.31 ;
      RECT  11.16 1.31 11.875 1.315 ;
      RECT  11.155 1.315 11.875 1.32 ;
      RECT  11.15 1.32 11.875 1.325 ;
      RECT  11.145 1.325 11.875 1.33 ;
      RECT  11.14 1.33 11.875 1.335 ;
      RECT  11.135 1.335 11.875 1.34 ;
      RECT  11.13 1.34 11.875 1.345 ;
      RECT  11.125 1.345 11.875 1.35 ;
      RECT  5.99 0.37 6.33 0.445 ;
      RECT  5.99 0.445 10.195 0.675 ;
      RECT  9.965 0.675 10.195 1.35 ;
      RECT  9.965 1.35 11.875 1.52 ;
      RECT  9.965 1.52 11.275 1.525 ;
      RECT  9.965 1.525 11.27 1.53 ;
      RECT  9.965 1.53 11.265 1.535 ;
      RECT  9.965 1.535 11.26 1.54 ;
      RECT  9.965 1.54 11.255 1.545 ;
      RECT  9.965 1.545 11.25 1.55 ;
      RECT  9.965 1.55 11.245 1.555 ;
      RECT  9.965 1.555 11.24 1.56 ;
      RECT  9.965 1.56 11.235 1.565 ;
      RECT  9.965 1.565 11.23 1.57 ;
      RECT  9.965 1.57 11.225 1.575 ;
      RECT  9.965 1.575 11.22 1.58 ;
      RECT  13.325 0.37 14.17 0.6 ;
      RECT  13.325 0.6 13.555 1.29 ;
      RECT  12.205 1.29 13.555 1.52 ;
      RECT  12.205 1.52 12.435 1.93 ;
      RECT  9.14 1.75 9.48 1.93 ;
      RECT  8.285 1.93 12.435 2.16 ;
      RECT  11.38 1.75 11.72 1.93 ;
      RECT  8.285 2.16 8.515 2.69 ;
      RECT  9.965 2.16 10.195 3.5 ;
      RECT  14.95 0.37 15.29 0.6 ;
      RECT  14.95 0.6 15.18 1.005 ;
      RECT  14.445 1.005 15.18 1.235 ;
      RECT  14.445 1.235 14.675 1.75 ;
      RECT  13.62 1.75 14.675 1.98 ;
      RECT  13.885 1.98 14.115 3.245 ;
      RECT  13.62 3.245 14.115 3.475 ;
      RECT  2.42 1.005 5.0 1.235 ;
      RECT  3.96 1.47 8.78 1.7 ;
      RECT  1.68 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
      RECT  3.245 1.51 3.475 1.93 ;
      RECT  3.245 1.93 7.955 2.16 ;
      RECT  7.725 2.16 7.955 3.245 ;
      RECT  3.245 2.16 3.475 3.405 ;
      RECT  6.9 3.245 9.635 3.475 ;
      RECT  9.405 2.39 9.635 3.245 ;
      RECT  12.765 1.75 13.26 1.98 ;
      RECT  12.765 1.98 12.995 2.445 ;
      RECT  11.59 2.445 12.995 2.675 ;
      RECT  12.765 2.675 12.995 3.245 ;
      RECT  12.765 3.245 13.26 3.475 ;
      RECT  5.99 2.405 7.45 2.635 ;
      RECT  3.96 3.805 5.0 4.035 ;
      RECT  2.42 4.365 8.78 4.595 ;
      RECT  10.68 4.365 11.72 4.595 ;
      RECT  1.51 4.925 4.09 5.155 ;
      RECT  1.51 5.155 1.85 5.23 ;
      RECT  3.75 5.155 4.09 5.23 ;
  END
END MDN_LDNRBSBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_LDNRBSBQ_2
#      Description : D-latch, neg-gate, lo-async-clear, lo-async-set, q-only
#      Equation    : iq,iqn=latch(enable=!G,data_in=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDNRBSBQ_2
  CLASS CORE ;
  FOREIGN MDN_LDNRBSBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.87 2.445 5.21 2.66 ;
      RECT  4.87 2.66 5.715 2.675 ;
      RECT  4.925 2.675 5.715 2.94 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.62 1.565 15.5 1.795 ;
      RECT  14.445 1.795 14.675 3.245 ;
      RECT  13.62 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.565 0.37 7.45 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  0.39 0.37 0.73 0.6 ;
      RECT  0.42 0.6 0.7 1.005 ;
      RECT  0.42 1.005 1.795 1.235 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  9.14 4.365 9.635 4.595 ;
      RECT  9.405 4.595 9.635 5.46 ;
      RECT  9.405 5.46 12.435 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  10.525 -0.14 11.2 0.14 ;
      RECT  10.525 0.14 10.755 1.005 ;
      RECT  10.525 1.005 11.02 1.235 ;
      RECT  7.28 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 1.005 ;
      RECT  6.2 1.005 7.955 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  12.7 0.37 13.05 0.6 ;
      RECT  12.7 0.6 12.93 1.005 ;
      RECT  11.34 1.005 12.93 1.235 ;
      RECT  11.34 1.235 11.57 1.565 ;
      RECT  8.23 0.37 9.33 0.6 ;
      RECT  9.1 0.6 9.33 1.565 ;
      RECT  9.1 1.565 11.57 1.795 ;
      RECT  9.965 1.795 10.195 3.53 ;
      RECT  14.95 0.37 15.29 0.6 ;
      RECT  14.95 0.6 15.18 1.005 ;
      RECT  13.83 0.37 14.17 0.6 ;
      RECT  13.94 0.6 14.17 1.005 ;
      RECT  13.16 1.005 15.18 1.235 ;
      RECT  13.16 1.235 13.39 1.565 ;
      RECT  12.765 1.565 13.39 1.795 ;
      RECT  12.765 1.795 12.995 3.245 ;
      RECT  12.765 3.245 13.26 3.475 ;
      RECT  2.42 1.005 5.0 1.235 ;
      RECT  3.96 1.525 8.78 1.755 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
      RECT  3.245 1.51 3.475 1.985 ;
      RECT  3.245 1.985 7.955 2.215 ;
      RECT  7.725 2.215 7.955 2.405 ;
      RECT  3.245 2.215 3.475 3.53 ;
      RECT  7.725 2.405 9.69 2.635 ;
      RECT  7.725 2.635 7.955 3.245 ;
      RECT  6.9 3.245 7.955 3.475 ;
      RECT  3.96 3.245 5.0 3.475 ;
      RECT  1.565 3.805 10.195 4.035 ;
      RECT  1.565 4.035 1.795 4.365 ;
      RECT  9.965 4.035 10.195 4.925 ;
      RECT  0.18 1.565 0.675 1.795 ;
      RECT  0.445 1.795 0.675 4.365 ;
      RECT  0.18 4.365 1.795 4.595 ;
      RECT  9.965 4.925 11.93 5.155 ;
      RECT  11.59 5.155 11.93 5.23 ;
      RECT  2.42 4.365 8.78 4.595 ;
      RECT  10.68 4.365 11.72 4.595 ;
      RECT  1.51 4.925 4.09 5.155 ;
      RECT  1.51 5.155 1.85 5.23 ;
      RECT  3.75 5.155 4.09 5.23 ;
  END
END MDN_LDNRBSBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_LDNRBSBQ_4
#      Description : D-latch, neg-gate, lo-async-clear, lo-async-set, q-only
#      Equation    : iq,iqn=latch(enable=!G,data_in=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDNRBSBQ_4
  CLASS CORE ;
  FOREIGN MDN_LDNRBSBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.87 2.445 5.21 2.66 ;
      RECT  4.87 2.66 5.715 2.675 ;
      RECT  4.925 2.675 5.715 2.94 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.62 1.565 17.74 1.795 ;
      RECT  15.565 1.795 15.795 3.245 ;
      RECT  13.62 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.565 0.37 7.45 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  0.39 0.37 0.73 0.6 ;
      RECT  0.42 0.6 0.7 1.005 ;
      RECT  0.42 1.005 1.795 1.235 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  9.14 4.365 9.635 4.595 ;
      RECT  9.405 4.595 9.635 5.46 ;
      RECT  9.405 5.46 12.435 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  10.525 -0.14 11.2 0.14 ;
      RECT  10.525 0.14 10.755 0.89 ;
      RECT  10.525 0.89 11.02 1.11 ;
      RECT  10.68 1.11 11.02 1.12 ;
      RECT  7.28 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 1.005 ;
      RECT  6.2 1.005 7.955 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  11.34 1.005 12.94 1.235 ;
      RECT  11.34 1.235 11.57 1.565 ;
      RECT  8.23 0.37 9.33 0.6 ;
      RECT  9.1 0.6 9.33 1.565 ;
      RECT  9.1 1.565 11.57 1.795 ;
      RECT  9.965 1.795 10.195 3.53 ;
      RECT  14.95 0.37 16.41 0.6 ;
      RECT  2.42 1.005 5.0 1.235 ;
      RECT  3.96 1.525 8.78 1.755 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
      RECT  12.765 1.565 13.26 1.795 ;
      RECT  12.765 1.795 12.995 2.405 ;
      RECT  12.765 2.405 15.29 2.635 ;
      RECT  12.765 2.635 12.995 3.245 ;
      RECT  12.765 3.245 13.26 3.475 ;
      RECT  3.245 1.51 3.475 1.985 ;
      RECT  3.245 1.985 7.955 2.215 ;
      RECT  7.725 2.215 7.955 2.405 ;
      RECT  3.245 2.215 3.475 3.53 ;
      RECT  7.725 2.405 9.69 2.635 ;
      RECT  7.725 2.635 7.955 3.245 ;
      RECT  6.9 3.245 7.955 3.475 ;
      RECT  16.07 2.405 17.53 2.635 ;
      RECT  3.96 3.245 5.0 3.475 ;
      RECT  1.565 3.805 10.195 4.035 ;
      RECT  1.565 4.035 1.795 4.365 ;
      RECT  9.965 4.035 10.195 4.925 ;
      RECT  0.18 1.565 0.675 1.795 ;
      RECT  0.445 1.795 0.675 4.365 ;
      RECT  0.18 4.365 1.795 4.595 ;
      RECT  9.965 4.925 11.93 5.155 ;
      RECT  11.59 5.155 11.93 5.23 ;
      RECT  2.42 4.365 8.78 4.595 ;
      RECT  10.68 4.365 11.72 4.595 ;
      RECT  1.51 4.925 4.09 5.155 ;
      RECT  1.51 5.155 1.85 5.23 ;
      RECT  3.75 5.155 4.09 5.23 ;
  END
END MDN_LDNRBSBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_LDNSBQ_1
#      Description : D-latch, neg-gate, lo-async-set, q-only
#      Equation    : iq,iqn=latch(enable=!G,data_in=D,preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDNSBQ_1
  CLASS CORE ;
  FOREIGN MDN_LDNSBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.14 1.565 10.195 1.795 ;
      RECT  9.965 1.795 10.195 3.245 ;
      RECT  9.14 3.245 10.195 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  6.16 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  6.255 0.14 6.485 1.29 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 4.09 0.6 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  4.015 1.005 6.025 1.235 ;
      RECT  5.795 1.235 6.025 1.565 ;
      RECT  4.015 1.235 4.245 1.85 ;
      RECT  5.795 1.565 7.185 1.795 ;
      RECT  6.955 0.95 7.185 1.565 ;
      RECT  8.44 1.005 8.805 1.235 ;
      RECT  8.575 1.235 8.805 2.405 ;
      RECT  8.575 2.405 9.69 2.635 ;
      RECT  8.575 2.635 8.805 3.245 ;
      RECT  8.44 3.245 8.805 3.475 ;
      RECT  1.72 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 2.405 ;
      RECT  2.125 2.405 2.845 2.635 ;
      RECT  2.125 2.635 2.355 3.805 ;
      RECT  1.72 3.805 2.355 4.035 ;
      RECT  3.245 1.51 3.475 2.405 ;
      RECT  3.245 2.405 5.055 2.635 ;
      RECT  3.245 2.635 3.475 3.53 ;
      RECT  7.105 2.405 8.345 2.635 ;
      RECT  7.725 2.635 7.955 3.805 ;
      RECT  4.715 1.51 4.945 1.945 ;
      RECT  4.715 1.945 5.535 2.175 ;
      RECT  5.305 2.175 5.535 3.245 ;
      RECT  4.66 3.245 5.715 3.475 ;
      RECT  5.485 3.475 5.715 3.805 ;
      RECT  5.485 3.805 7.955 4.035 ;
      RECT  3.245 3.805 5.155 4.035 ;
      RECT  3.245 4.035 3.475 4.365 ;
      RECT  4.925 4.035 5.155 4.365 ;
      RECT  2.42 4.365 3.475 4.595 ;
      RECT  4.925 4.365 7.24 4.595 ;
      RECT  0.18 4.365 1.795 4.595 ;
      RECT  1.565 4.595 1.795 4.925 ;
      RECT  1.565 4.925 4.245 5.155 ;
      RECT  4.015 4.31 4.245 4.925 ;
  END
END MDN_LDNSBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_LDNSBQ_2
#      Description : D-latch, neg-gate, lo-async-set, q-only
#      Equation    : iq,iqn=latch(enable=!G,data_in=D,preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDNSBQ_2
  CLASS CORE ;
  FOREIGN MDN_LDNSBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.14 1.565 11.02 1.795 ;
      RECT  9.405 1.795 9.635 3.245 ;
      RECT  9.14 3.245 11.02 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  4.66 4.365 6.54 4.595 ;
      RECT  4.925 4.595 5.155 5.46 ;
      RECT  4.925 5.46 7.955 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.735 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  6.16 -0.14 7.28 0.14 ;
      RECT  6.255 0.14 6.485 1.29 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.445 ;
      RECT  1.51 0.445 4.09 0.675 ;
      RECT  3.75 0.37 4.09 0.445 ;
      RECT  10.47 0.37 10.81 0.6 ;
      RECT  10.525 0.6 10.755 1.005 ;
      RECT  9.35 0.37 9.69 0.6 ;
      RECT  9.405 0.6 9.635 1.005 ;
      RECT  8.285 1.005 10.755 1.235 ;
      RECT  8.285 1.235 8.515 3.245 ;
      RECT  8.285 3.245 8.78 3.475 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.005 6.01 1.235 ;
      RECT  5.78 1.235 6.01 1.565 ;
      RECT  5.78 1.565 7.24 1.795 ;
      RECT  1.715 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.805 ;
      RECT  1.72 3.805 2.915 4.035 ;
      RECT  4.66 1.565 5.55 1.795 ;
      RECT  5.32 1.795 5.55 2.125 ;
      RECT  5.32 2.125 5.715 2.355 ;
      RECT  5.485 2.355 5.715 3.53 ;
      RECT  3.245 1.51 3.475 2.405 ;
      RECT  3.245 2.405 5.08 2.635 ;
      RECT  3.245 2.635 3.475 3.53 ;
      RECT  3.245 3.805 7.24 4.035 ;
      RECT  3.245 4.035 3.475 4.365 ;
      RECT  2.42 4.365 3.475 4.595 ;
      RECT  0.18 4.365 1.795 4.595 ;
      RECT  1.565 4.595 1.795 4.925 ;
      RECT  1.565 4.925 4.245 5.155 ;
      RECT  4.015 4.31 4.245 4.925 ;
      RECT  7.22 4.365 8.515 4.595 ;
      RECT  7.22 4.595 7.45 5.0 ;
      RECT  8.285 4.595 8.515 5.0 ;
      RECT  5.425 5.0 7.45 5.23 ;
      RECT  8.23 5.0 8.57 5.23 ;
  END
END MDN_LDNSBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_LDNSBQ_4
#      Description : D-latch, neg-gate, lo-async-set, q-only
#      Equation    : iq,iqn=latch(enable=!G,data_in=D,preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDNSBQ_4
  CLASS CORE ;
  FOREIGN MDN_LDNSBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.14 1.565 13.265 1.795 ;
      RECT  11.085 1.795 11.315 3.245 ;
      RECT  9.14 3.245 13.26 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  4.655 4.365 6.54 4.595 ;
      RECT  4.925 4.595 5.155 5.46 ;
      RECT  4.925 5.46 7.955 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  9.965 -0.14 11.2 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  6.16 -0.14 7.28 0.14 ;
      RECT  6.255 0.14 6.485 1.29 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 4.09 0.6 ;
      RECT  10.47 0.37 11.93 0.6 ;
      RECT  0.175 1.005 2.76 1.235 ;
      RECT  3.96 1.005 6.025 1.235 ;
      RECT  5.795 1.235 6.025 1.565 ;
      RECT  5.795 1.565 7.24 1.795 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.805 ;
      RECT  1.72 3.805 2.915 4.035 ;
      RECT  4.66 1.565 5.565 1.795 ;
      RECT  5.335 1.795 5.565 2.125 ;
      RECT  5.335 2.125 5.715 2.355 ;
      RECT  5.485 2.355 5.715 3.53 ;
      RECT  8.285 1.565 8.78 1.795 ;
      RECT  8.285 1.795 8.515 2.405 ;
      RECT  8.285 2.405 10.65 2.635 ;
      RECT  8.285 2.635 8.515 3.245 ;
      RECT  8.285 3.245 8.78 3.475 ;
      RECT  3.245 1.51 3.475 2.405 ;
      RECT  3.245 2.405 5.07 2.635 ;
      RECT  3.245 2.635 3.475 3.53 ;
      RECT  11.7 2.405 13.05 2.635 ;
      RECT  3.245 3.805 7.24 4.035 ;
      RECT  3.245 4.035 3.475 4.365 ;
      RECT  2.42 4.365 3.475 4.595 ;
      RECT  0.18 4.365 1.795 4.595 ;
      RECT  1.565 4.595 1.795 4.925 ;
      RECT  1.565 4.925 4.245 5.155 ;
      RECT  4.015 4.31 4.245 4.925 ;
      RECT  7.22 4.365 8.46 4.595 ;
      RECT  7.22 4.595 7.45 5.0 ;
      RECT  8.23 4.595 8.46 5.0 ;
      RECT  5.43 5.0 7.45 5.23 ;
      RECT  8.23 5.0 8.57 5.23 ;
  END
END MDN_LDNSBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_LDPQ_4
#      Description : D-latch, pos-gate, q-only
#      Equation    : iq,iqn=latch(enable=G,data_in=D):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDPQ_4
  CLASS CORE ;
  FOREIGN MDN_LDPQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.44 1.565 11.72 1.795 ;
      RECT  11.085 1.795 11.315 3.245 ;
      RECT  8.44 3.245 11.72 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 2.97 0.6 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.005 6.54 1.235 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 2.685 ;
      RECT  2.685 2.685 3.97 2.915 ;
      RECT  3.74 2.345 3.97 2.685 ;
      RECT  2.685 2.915 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
      RECT  3.19 1.565 4.43 1.795 ;
      RECT  4.2 1.795 4.43 2.405 ;
      RECT  4.2 2.405 5.21 2.635 ;
      RECT  4.2 2.635 4.43 3.245 ;
      RECT  3.19 3.245 4.43 3.475 ;
      RECT  4.66 1.565 6.275 1.795 ;
      RECT  6.045 1.795 6.275 3.245 ;
      RECT  4.66 3.245 6.275 3.475 ;
      RECT  6.955 1.51 7.185 2.685 ;
      RECT  6.955 2.685 10.755 2.915 ;
      RECT  8.285 2.35 8.515 2.685 ;
      RECT  9.405 2.35 9.635 2.685 ;
      RECT  10.525 2.35 10.755 2.685 ;
      RECT  6.955 2.915 7.185 3.53 ;
      RECT  2.42 3.805 6.54 4.035 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  5.99 5.0 7.45 5.23 ;
      RECT  10.47 5.0 11.93 5.23 ;
  END
END MDN_LDPQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_LDPQ_1
#      Description : D-latch, pos-gate, q-only
#      Equation    : iq,iqn=latch(enable=G,data_in=D):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDPQ_1
  CLASS CORE ;
  FOREIGN MDN_LDPQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.605 1.565 7.24 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  6.605 3.245 7.24 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  8.4 5.46 9.13 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 2.97 0.6 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.005 6.54 1.235 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 2.685 ;
      RECT  2.685 2.685 3.97 2.915 ;
      RECT  3.74 2.35 3.97 2.685 ;
      RECT  2.685 2.915 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
      RECT  3.19 1.565 4.43 1.795 ;
      RECT  4.2 1.795 4.43 2.685 ;
      RECT  4.2 2.685 5.155 2.915 ;
      RECT  4.925 2.35 5.155 2.685 ;
      RECT  4.2 2.915 4.43 3.245 ;
      RECT  3.19 3.245 4.43 3.475 ;
      RECT  4.66 1.565 5.715 1.795 ;
      RECT  5.485 1.795 5.715 2.405 ;
      RECT  5.485 2.405 6.33 2.635 ;
      RECT  5.485 2.635 5.715 3.245 ;
      RECT  4.66 3.245 5.715 3.475 ;
      RECT  2.42 3.805 6.54 4.035 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.925 4.365 6.275 4.595 ;
      RECT  4.925 4.595 5.155 4.925 ;
      RECT  6.045 4.595 6.275 5.0 ;
      RECT  3.19 4.925 5.155 5.155 ;
      RECT  6.045 5.0 7.45 5.23 ;
  END
END MDN_LDPQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_LDPQ_2
#      Description : D-latch, pos-gate, q-only
#      Equation    : iq,iqn=latch(enable=G,data_in=D):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDPQ_2
  CLASS CORE ;
  FOREIGN MDN_LDPQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 8.78 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  6.9 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  8.4 5.46 9.13 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 2.97 0.6 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.005 6.54 1.235 ;
      RECT  1.72 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 2.685 ;
      RECT  2.125 2.685 3.97 2.915 ;
      RECT  3.74 2.35 3.97 2.685 ;
      RECT  2.125 2.915 2.355 3.245 ;
      RECT  1.72 3.245 2.355 3.475 ;
      RECT  3.19 1.565 4.43 1.795 ;
      RECT  4.2 1.795 4.43 2.405 ;
      RECT  4.2 2.405 5.21 2.635 ;
      RECT  4.2 2.635 4.43 3.245 ;
      RECT  3.19 3.245 4.43 3.475 ;
      RECT  4.66 1.565 6.275 1.795 ;
      RECT  6.045 1.795 6.275 3.245 ;
      RECT  4.66 3.245 6.275 3.475 ;
      RECT  2.42 3.805 6.54 4.035 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.98 4.365 8.46 4.595 ;
      RECT  4.98 4.595 5.21 5.0 ;
      RECT  7.22 4.595 7.45 5.0 ;
      RECT  8.23 4.595 8.46 5.0 ;
      RECT  4.87 5.0 5.21 5.23 ;
      RECT  7.11 5.0 7.45 5.23 ;
      RECT  8.23 5.0 8.57 5.23 ;
  END
END MDN_LDPQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_LDPRBQ_4
#      Description : D-latch, pos-gate, lo-async-clear, q-only
#      Equation    : iq,iqn=latch(enable=G,data_in=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDPRBQ_4
  CLASS CORE ;
  FOREIGN MDN_LDPRBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 7.42 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.38 1.565 15.5 1.795 ;
      RECT  13.325 1.795 13.555 3.245 ;
      RECT  11.38 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.605 0.37 8.57 0.6 ;
      RECT  6.605 0.6 6.835 1.005 ;
      RECT  3.245 1.005 6.835 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  2.66 1.565 3.475 1.795 ;
      RECT  2.66 1.795 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  6.55 5.46 7.955 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  8.4 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  8.845 0.14 9.075 1.005 ;
      RECT  8.44 1.005 9.075 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 1.005 ;
      RECT  1.005 1.005 2.76 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.445 ;
      RECT  1.51 0.445 6.33 0.675 ;
      RECT  5.99 0.37 6.33 0.445 ;
      RECT  10.47 0.37 10.81 0.6 ;
      RECT  10.47 0.6 10.7 1.005 ;
      RECT  9.405 1.005 10.7 1.235 ;
      RECT  9.405 1.235 9.635 1.565 ;
      RECT  8.285 1.565 9.635 1.795 ;
      RECT  8.285 1.795 8.515 3.245 ;
      RECT  9.405 1.795 9.635 3.245 ;
      RECT  6.045 3.245 8.515 3.475 ;
      RECT  9.14 3.245 9.635 3.475 ;
      RECT  6.045 3.475 6.275 3.49 ;
      RECT  3.805 2.35 4.035 3.49 ;
      RECT  3.805 3.49 6.275 3.72 ;
      RECT  12.71 0.37 14.17 0.6 ;
      RECT  1.72 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 4.41 ;
      RECT  1.72 4.41 4.03 4.64 ;
      RECT  3.8 4.64 4.03 4.925 ;
      RECT  3.8 4.925 5.2 5.155 ;
      RECT  4.86 5.155 5.2 5.23 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  10.735 1.51 10.965 2.125 ;
      RECT  10.735 2.125 12.995 2.355 ;
      RECT  11.645 2.355 11.875 2.69 ;
      RECT  12.765 2.355 12.995 2.69 ;
      RECT  10.735 2.355 10.965 3.53 ;
      RECT  13.885 2.125 15.235 2.355 ;
      RECT  13.885 2.355 14.115 2.69 ;
      RECT  15.005 2.355 15.235 2.69 ;
      RECT  5.485 1.51 5.715 3.03 ;
      RECT  5.43 3.03 5.77 3.26 ;
      RECT  6.795 3.805 7.24 4.035 ;
      RECT  6.795 4.035 7.025 4.41 ;
      RECT  4.66 4.41 7.025 4.64 ;
      RECT  3.96 3.95 6.54 4.18 ;
      RECT  7.255 4.365 9.075 4.595 ;
      RECT  7.255 4.595 7.485 5.0 ;
      RECT  8.845 4.595 9.075 5.0 ;
      RECT  5.43 5.0 7.485 5.23 ;
      RECT  8.845 5.0 9.69 5.23 ;
  END
END MDN_LDPRBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_LDPRBQ_1
#      Description : D-latch, pos-gate, lo-async-clear, q-only
#      Equation    : iq,iqn=latch(enable=G,data_in=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDPRBQ_1
  CLASS CORE ;
  FOREIGN MDN_LDPRBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 7.42 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.525 1.565 11.02 1.795 ;
      RECT  10.525 1.795 10.755 3.245 ;
      RECT  10.525 3.245 11.02 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.605 0.37 8.57 0.6 ;
      RECT  6.605 0.6 6.835 1.005 ;
      RECT  3.245 1.005 6.835 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  2.685 1.565 3.475 1.795 ;
      RECT  2.685 1.795 2.915 2.125 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  6.55 5.46 7.955 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  8.4 -0.14 9.52 0.14 ;
      RECT  8.845 0.14 9.075 1.005 ;
      RECT  8.44 1.005 9.075 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 1.005 ;
      RECT  1.005 1.005 2.76 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.445 ;
      RECT  1.51 0.445 6.33 0.675 ;
      RECT  5.99 0.37 6.33 0.445 ;
      RECT  1.72 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 4.41 ;
      RECT  1.72 4.41 4.035 4.64 ;
      RECT  3.805 4.64 4.035 4.925 ;
      RECT  3.805 4.925 5.2 5.155 ;
      RECT  4.86 5.155 5.2 5.23 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  9.14 1.565 9.635 1.795 ;
      RECT  9.405 1.795 9.635 3.805 ;
      RECT  6.045 3.245 7.955 3.475 ;
      RECT  6.045 3.475 6.275 3.49 ;
      RECT  7.725 3.475 7.955 3.805 ;
      RECT  3.805 2.35 4.035 3.49 ;
      RECT  3.805 3.49 6.275 3.72 ;
      RECT  7.725 3.805 9.635 4.035 ;
      RECT  5.485 1.51 5.715 3.03 ;
      RECT  5.43 3.03 5.77 3.26 ;
      RECT  6.795 3.805 7.24 4.035 ;
      RECT  6.795 4.035 7.025 4.41 ;
      RECT  4.66 4.41 7.025 4.64 ;
      RECT  3.96 3.95 6.54 4.18 ;
      RECT  7.255 4.365 10.7 4.595 ;
      RECT  7.255 4.595 7.485 4.925 ;
      RECT  9.46 4.595 9.69 5.0 ;
      RECT  10.47 4.595 10.7 5.0 ;
      RECT  5.43 4.925 7.485 5.155 ;
      RECT  9.35 5.0 9.69 5.23 ;
      RECT  10.47 5.0 10.81 5.23 ;
  END
END MDN_LDPRBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_LDPRBQ_2
#      Description : D-latch, pos-gate, lo-async-clear, q-only
#      Equation    : iq,iqn=latch(enable=G,data_in=D,clear=!RD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDPRBQ_2
  CLASS CORE ;
  FOREIGN MDN_LDPRBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.925 2.125 6.3 2.355 ;
      RECT  4.925 2.355 5.155 2.69 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.11 0.37 7.45 0.6 ;
      RECT  7.14 0.6 7.42 1.235 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.14 1.565 11.02 1.795 ;
      RECT  9.965 1.795 10.195 3.245 ;
      RECT  9.14 3.245 11.02 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  5.79 0.37 6.33 0.445 ;
      RECT  1.005 0.445 6.33 0.675 ;
      RECT  1.005 0.675 1.235 1.565 ;
      RECT  0.415 1.565 1.235 1.795 ;
      RECT  0.42 1.795 0.7 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.43 5.135 5.77 5.46 ;
      RECT  5.04 5.46 6.16 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  6.55 -0.14 7.28 0.14 ;
      RECT  6.605 0.14 6.835 1.005 ;
      RECT  6.2 1.005 6.835 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  3.32 1.005 5.715 1.01 ;
      RECT  3.315 1.01 5.715 1.015 ;
      RECT  3.31 1.015 5.715 1.02 ;
      RECT  3.305 1.02 5.715 1.025 ;
      RECT  3.3 1.025 5.715 1.03 ;
      RECT  3.295 1.03 5.715 1.035 ;
      RECT  3.29 1.035 5.715 1.04 ;
      RECT  3.285 1.04 5.715 1.045 ;
      RECT  3.28 1.045 5.715 1.05 ;
      RECT  3.275 1.05 5.715 1.055 ;
      RECT  3.27 1.055 5.715 1.06 ;
      RECT  3.265 1.06 5.715 1.065 ;
      RECT  3.26 1.065 5.715 1.07 ;
      RECT  3.255 1.07 5.715 1.075 ;
      RECT  3.25 1.075 5.715 1.08 ;
      RECT  3.245 1.08 5.715 1.085 ;
      RECT  3.24 1.085 5.715 1.09 ;
      RECT  3.235 1.09 5.715 1.095 ;
      RECT  3.23 1.095 5.715 1.1 ;
      RECT  3.225 1.1 5.715 1.105 ;
      RECT  3.22 1.105 5.715 1.11 ;
      RECT  3.215 1.11 5.715 1.115 ;
      RECT  3.21 1.115 5.715 1.12 ;
      RECT  3.205 1.12 5.715 1.125 ;
      RECT  3.2 1.125 5.715 1.13 ;
      RECT  3.195 1.13 5.715 1.135 ;
      RECT  3.19 1.135 5.715 1.14 ;
      RECT  3.185 1.14 5.715 1.145 ;
      RECT  3.18 1.145 5.715 1.15 ;
      RECT  3.175 1.15 5.715 1.155 ;
      RECT  3.17 1.155 5.715 1.16 ;
      RECT  3.165 1.16 5.715 1.165 ;
      RECT  3.16 1.165 5.715 1.17 ;
      RECT  3.155 1.17 5.715 1.175 ;
      RECT  3.15 1.175 5.715 1.18 ;
      RECT  3.145 1.18 5.715 1.185 ;
      RECT  3.14 1.185 5.715 1.19 ;
      RECT  3.135 1.19 5.715 1.195 ;
      RECT  3.13 1.195 5.715 1.2 ;
      RECT  3.125 1.2 5.715 1.205 ;
      RECT  3.12 1.205 5.715 1.21 ;
      RECT  3.115 1.21 5.715 1.215 ;
      RECT  3.11 1.215 5.715 1.22 ;
      RECT  3.105 1.22 5.715 1.225 ;
      RECT  3.1 1.225 5.715 1.23 ;
      RECT  3.095 1.23 5.715 1.235 ;
      RECT  3.09 1.235 3.415 1.24 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  3.085 1.24 3.41 1.245 ;
      RECT  3.08 1.245 3.405 1.25 ;
      RECT  3.075 1.25 3.4 1.255 ;
      RECT  3.07 1.255 3.395 1.26 ;
      RECT  3.065 1.26 3.39 1.265 ;
      RECT  3.06 1.265 3.385 1.27 ;
      RECT  3.055 1.27 3.38 1.275 ;
      RECT  3.05 1.275 3.375 1.28 ;
      RECT  3.045 1.28 3.37 1.285 ;
      RECT  3.04 1.285 3.365 1.29 ;
      RECT  3.035 1.29 3.36 1.295 ;
      RECT  3.03 1.295 3.355 1.3 ;
      RECT  3.025 1.3 3.35 1.305 ;
      RECT  3.02 1.305 3.345 1.31 ;
      RECT  3.015 1.31 3.34 1.315 ;
      RECT  3.01 1.315 3.335 1.32 ;
      RECT  3.005 1.32 3.33 1.325 ;
      RECT  3.0 1.325 3.325 1.33 ;
      RECT  2.995 1.33 3.32 1.335 ;
      RECT  2.99 1.335 3.315 1.34 ;
      RECT  2.985 1.34 3.31 1.345 ;
      RECT  2.98 1.345 3.305 1.35 ;
      RECT  2.975 1.35 3.3 1.355 ;
      RECT  2.97 1.355 3.295 1.36 ;
      RECT  2.965 1.36 3.29 1.365 ;
      RECT  2.96 1.365 3.285 1.37 ;
      RECT  2.955 1.37 3.28 1.375 ;
      RECT  2.95 1.375 3.275 1.38 ;
      RECT  2.945 1.38 3.27 1.385 ;
      RECT  2.94 1.385 3.265 1.39 ;
      RECT  2.935 1.39 3.26 1.395 ;
      RECT  2.93 1.395 3.255 1.4 ;
      RECT  2.925 1.4 3.25 1.405 ;
      RECT  2.92 1.405 3.245 1.41 ;
      RECT  2.915 1.41 3.24 1.415 ;
      RECT  2.91 1.415 3.235 1.42 ;
      RECT  2.905 1.42 3.23 1.425 ;
      RECT  2.9 1.425 3.225 1.43 ;
      RECT  2.895 1.43 3.22 1.435 ;
      RECT  2.89 1.435 3.215 1.44 ;
      RECT  2.885 1.44 3.21 1.445 ;
      RECT  2.88 1.445 3.205 1.45 ;
      RECT  2.875 1.45 3.2 1.455 ;
      RECT  2.87 1.455 3.195 1.46 ;
      RECT  2.865 1.46 3.19 1.465 ;
      RECT  2.86 1.465 3.185 1.47 ;
      RECT  2.855 1.47 3.18 1.475 ;
      RECT  2.85 1.475 3.175 1.48 ;
      RECT  2.845 1.48 3.17 1.485 ;
      RECT  2.84 1.485 3.165 1.49 ;
      RECT  2.835 1.49 3.16 1.495 ;
      RECT  2.83 1.495 3.155 1.5 ;
      RECT  2.825 1.5 3.15 1.505 ;
      RECT  2.82 1.505 3.145 1.51 ;
      RECT  2.815 1.51 3.14 1.515 ;
      RECT  2.81 1.515 3.135 1.52 ;
      RECT  2.805 1.52 3.13 1.525 ;
      RECT  2.8 1.525 3.125 1.53 ;
      RECT  2.795 1.53 3.12 1.535 ;
      RECT  2.79 1.535 3.115 1.54 ;
      RECT  2.785 1.54 3.11 1.545 ;
      RECT  2.78 1.545 3.105 1.55 ;
      RECT  2.775 1.55 3.1 1.555 ;
      RECT  2.77 1.555 3.095 1.56 ;
      RECT  2.765 1.56 3.09 1.565 ;
      RECT  2.76 1.565 3.085 1.57 ;
      RECT  5.485 1.565 7.395 1.795 ;
      RECT  2.755 1.57 3.08 1.575 ;
      RECT  2.75 1.575 3.075 1.58 ;
      RECT  2.745 1.58 3.07 1.585 ;
      RECT  2.74 1.585 3.065 1.59 ;
      RECT  2.735 1.59 3.06 1.595 ;
      RECT  2.73 1.595 3.055 1.6 ;
      RECT  2.725 1.6 3.05 1.605 ;
      RECT  2.72 1.605 3.045 1.61 ;
      RECT  2.715 1.61 3.04 1.615 ;
      RECT  2.71 1.615 3.035 1.62 ;
      RECT  2.705 1.62 3.03 1.625 ;
      RECT  2.7 1.625 3.025 1.63 ;
      RECT  2.695 1.63 3.02 1.635 ;
      RECT  2.69 1.635 3.015 1.64 ;
      RECT  2.685 1.64 3.01 1.645 ;
      RECT  2.685 1.645 3.005 1.65 ;
      RECT  2.685 1.65 3.0 1.655 ;
      RECT  2.685 1.655 2.995 1.66 ;
      RECT  2.685 1.66 2.99 1.665 ;
      RECT  2.685 1.665 2.985 1.67 ;
      RECT  2.685 1.67 2.98 1.675 ;
      RECT  2.685 1.675 2.975 1.68 ;
      RECT  2.685 1.68 2.97 1.685 ;
      RECT  2.685 1.685 2.965 1.69 ;
      RECT  2.685 1.69 2.96 1.695 ;
      RECT  2.685 1.695 2.955 1.7 ;
      RECT  2.685 1.7 2.95 1.705 ;
      RECT  2.685 1.705 2.945 1.71 ;
      RECT  2.685 1.71 2.94 1.715 ;
      RECT  2.685 1.715 2.935 1.72 ;
      RECT  2.685 1.72 2.93 1.725 ;
      RECT  2.685 1.725 2.925 1.73 ;
      RECT  2.685 1.73 2.92 1.735 ;
      RECT  2.685 1.735 2.915 2.695 ;
      RECT  7.165 1.795 7.395 3.245 ;
      RECT  6.9 3.245 7.395 3.475 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  8.285 1.565 8.78 1.795 ;
      RECT  8.285 1.795 8.515 3.245 ;
      RECT  8.285 3.245 8.78 3.475 ;
      RECT  3.295 1.695 3.525 3.03 ;
      RECT  3.19 3.03 5.715 3.26 ;
      RECT  5.485 3.26 5.715 3.755 ;
      RECT  5.485 3.755 9.69 3.985 ;
      RECT  9.46 3.985 9.69 4.365 ;
      RECT  9.46 4.365 10.7 4.595 ;
      RECT  9.46 4.595 9.69 5.0 ;
      RECT  10.47 4.595 10.7 5.0 ;
      RECT  8.23 5.0 9.69 5.23 ;
      RECT  10.47 5.0 10.81 5.23 ;
      RECT  2.42 3.49 5.0 3.72 ;
      RECT  2.685 3.95 4.245 4.18 ;
      RECT  4.015 4.18 4.245 4.29 ;
      RECT  2.685 4.18 2.915 4.365 ;
      RECT  1.72 4.365 2.915 4.595 ;
      RECT  4.51 4.215 8.78 4.445 ;
      RECT  4.51 4.445 4.74 4.54 ;
      RECT  3.245 4.54 4.74 4.77 ;
      RECT  3.245 4.77 3.475 5.0 ;
      RECT  1.51 5.0 3.475 5.23 ;
      RECT  4.97 4.675 6.275 4.905 ;
      RECT  4.97 4.905 5.2 5.0 ;
      RECT  6.045 4.905 6.275 5.0 ;
      RECT  3.75 5.0 5.2 5.23 ;
      RECT  6.045 5.0 7.45 5.23 ;
  END
END MDN_LDPRBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_LDPRBSBQ_1
#      Description : D-latch, pos-gate, lo-async-clear, lo-async-set, q-only
#      Equation    : iq,iqn=latch(enable=G,data_in=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDPRBSBQ_1
  CLASS CORE ;
  FOREIGN MDN_LDPRBSBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.925 2.39 5.155 2.685 ;
      RECT  4.925 2.685 5.74 2.915 ;
      RECT  5.46 2.915 5.74 3.475 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 3.245 ;
      RECT  15.005 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.74 4.365 13.02 5.0 ;
      RECT  12.71 5.0 13.05 5.23 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.39 10.78 3.475 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.14 4.365 9.635 4.595 ;
      RECT  9.405 4.595 9.635 5.46 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 9.635 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.205 -0.14 13.44 0.14 ;
      RECT  12.205 0.14 12.435 0.6 ;
      RECT  10.08 -0.14 10.755 0.14 ;
      RECT  10.525 0.14 10.755 0.89 ;
      RECT  10.525 0.89 11.02 1.12 ;
      RECT  5.6 -0.14 6.72 0.14 ;
      RECT  6.045 0.14 6.275 1.005 ;
      RECT  6.045 1.005 7.24 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.09 0.445 ;
      RECT  1.565 0.445 4.09 0.675 ;
      RECT  1.565 0.675 1.795 1.565 ;
      RECT  1.565 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 0.83 ;
      RECT  11.25 0.83 12.94 1.06 ;
      RECT  11.25 1.06 11.48 1.225 ;
      RECT  11.245 1.225 11.48 1.23 ;
      RECT  11.24 1.23 11.48 1.235 ;
      RECT  11.235 1.235 11.48 1.24 ;
      RECT  11.23 1.24 11.48 1.245 ;
      RECT  11.225 1.245 11.48 1.25 ;
      RECT  11.22 1.25 11.48 1.255 ;
      RECT  11.215 1.255 11.48 1.26 ;
      RECT  11.21 1.26 11.48 1.265 ;
      RECT  11.205 1.265 11.48 1.27 ;
      RECT  11.2 1.27 11.48 1.275 ;
      RECT  11.195 1.275 11.48 1.28 ;
      RECT  11.19 1.28 11.48 1.285 ;
      RECT  11.185 1.285 11.48 1.29 ;
      RECT  11.18 1.29 11.48 1.295 ;
      RECT  11.175 1.295 11.48 1.3 ;
      RECT  11.17 1.3 11.48 1.305 ;
      RECT  11.165 1.305 11.48 1.31 ;
      RECT  11.16 1.31 11.48 1.315 ;
      RECT  11.155 1.315 11.48 1.32 ;
      RECT  11.15 1.32 11.475 1.325 ;
      RECT  11.145 1.325 11.47 1.33 ;
      RECT  11.14 1.33 11.465 1.335 ;
      RECT  11.135 1.335 11.46 1.34 ;
      RECT  11.13 1.34 11.455 1.345 ;
      RECT  11.125 1.345 11.45 1.35 ;
      RECT  7.11 0.37 7.45 0.445 ;
      RECT  7.11 0.445 10.195 0.675 ;
      RECT  9.965 0.675 10.195 1.35 ;
      RECT  9.965 1.35 11.445 1.355 ;
      RECT  9.965 1.355 11.44 1.36 ;
      RECT  9.965 1.36 11.435 1.365 ;
      RECT  9.965 1.365 11.43 1.37 ;
      RECT  9.965 1.37 11.425 1.375 ;
      RECT  9.965 1.375 11.42 1.38 ;
      RECT  9.965 1.38 11.415 1.385 ;
      RECT  9.965 1.385 11.41 1.39 ;
      RECT  9.965 1.39 11.405 1.395 ;
      RECT  9.965 1.395 11.4 1.4 ;
      RECT  9.965 1.4 11.395 1.405 ;
      RECT  9.965 1.405 11.39 1.41 ;
      RECT  9.965 1.41 11.385 1.415 ;
      RECT  9.965 1.415 11.38 1.42 ;
      RECT  9.965 1.42 11.375 1.425 ;
      RECT  9.965 1.425 11.37 1.43 ;
      RECT  9.965 1.43 11.365 1.435 ;
      RECT  9.965 1.435 11.36 1.44 ;
      RECT  9.965 1.44 11.355 1.445 ;
      RECT  9.965 1.445 11.35 1.45 ;
      RECT  9.965 1.45 11.345 1.455 ;
      RECT  9.965 1.455 11.34 1.46 ;
      RECT  9.965 1.46 11.335 1.465 ;
      RECT  9.965 1.465 11.33 1.47 ;
      RECT  9.965 1.47 11.325 1.475 ;
      RECT  9.965 1.475 11.32 1.48 ;
      RECT  9.965 1.48 11.315 1.485 ;
      RECT  9.965 1.485 11.31 1.49 ;
      RECT  9.965 1.49 11.305 1.495 ;
      RECT  9.965 1.495 11.3 1.5 ;
      RECT  9.965 1.5 11.295 1.505 ;
      RECT  9.965 1.505 11.29 1.51 ;
      RECT  9.965 1.51 11.285 1.515 ;
      RECT  9.965 1.515 11.28 1.52 ;
      RECT  9.965 1.52 11.275 1.525 ;
      RECT  9.965 1.525 11.27 1.53 ;
      RECT  9.965 1.53 11.265 1.535 ;
      RECT  9.965 1.535 11.26 1.54 ;
      RECT  9.965 1.54 11.255 1.545 ;
      RECT  9.965 1.545 11.25 1.55 ;
      RECT  9.965 1.55 11.245 1.555 ;
      RECT  9.965 1.555 11.24 1.56 ;
      RECT  9.965 1.56 11.235 1.565 ;
      RECT  9.965 1.565 11.23 1.57 ;
      RECT  9.965 1.57 11.225 1.575 ;
      RECT  9.965 1.575 11.22 1.58 ;
      RECT  13.325 0.37 14.17 0.6 ;
      RECT  13.325 0.6 13.555 1.29 ;
      RECT  12.205 1.29 13.555 1.52 ;
      RECT  12.205 1.52 12.435 1.925 ;
      RECT  9.14 1.745 9.48 1.925 ;
      RECT  8.285 1.925 12.435 2.155 ;
      RECT  11.38 1.75 11.72 1.925 ;
      RECT  8.285 2.155 8.515 2.69 ;
      RECT  9.965 2.155 10.195 3.53 ;
      RECT  14.95 0.37 15.29 0.6 ;
      RECT  14.95 0.6 15.18 1.005 ;
      RECT  13.885 1.005 15.18 1.235 ;
      RECT  13.885 1.235 14.115 1.75 ;
      RECT  13.62 1.75 14.115 1.98 ;
      RECT  13.885 1.98 14.115 3.245 ;
      RECT  13.62 3.245 14.115 3.475 ;
      RECT  2.42 1.005 5.0 1.235 ;
      RECT  3.96 1.465 8.78 1.695 ;
      RECT  3.245 1.51 3.475 1.925 ;
      RECT  3.245 1.925 7.955 2.155 ;
      RECT  7.725 2.155 7.955 3.245 ;
      RECT  3.245 2.155 3.475 3.405 ;
      RECT  6.9 3.245 9.635 3.475 ;
      RECT  9.405 2.39 9.635 3.245 ;
      RECT  12.765 1.75 13.26 1.98 ;
      RECT  12.765 1.98 12.995 2.445 ;
      RECT  11.59 2.445 12.995 2.675 ;
      RECT  12.765 2.675 12.995 3.245 ;
      RECT  12.765 3.245 13.26 3.475 ;
      RECT  5.99 2.405 7.45 2.635 ;
      RECT  3.96 3.245 5.0 3.475 ;
      RECT  2.42 4.365 8.78 4.595 ;
      RECT  10.68 4.365 11.72 4.595 ;
      RECT  1.51 5.0 2.97 5.23 ;
  END
END MDN_LDPRBSBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_LDPRBSBQ_2
#      Description : D-latch, pos-gate, lo-async-clear, lo-async-set, q-only
#      Equation    : iq,iqn=latch(enable=G,data_in=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDPRBSBQ_2
  CLASS CORE ;
  FOREIGN MDN_LDPRBSBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.915 2.385 5.165 2.66 ;
      RECT  4.915 2.66 5.715 2.665 ;
      RECT  4.925 2.665 5.715 2.94 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.62 1.565 15.5 1.795 ;
      RECT  14.445 1.795 14.675 3.245 ;
      RECT  13.62 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.565 0.37 7.45 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  0.39 0.37 0.73 0.6 ;
      RECT  0.42 0.6 0.7 1.005 ;
      RECT  0.42 1.005 1.795 1.235 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  9.14 4.365 9.635 4.595 ;
      RECT  9.405 4.595 9.635 5.46 ;
      RECT  9.405 5.46 12.435 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  10.525 -0.14 11.2 0.14 ;
      RECT  10.525 0.14 10.755 1.005 ;
      RECT  10.525 1.005 11.02 1.235 ;
      RECT  7.28 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 1.005 ;
      RECT  6.2 1.005 7.955 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  12.7 0.37 13.05 0.6 ;
      RECT  12.7 0.6 12.93 1.005 ;
      RECT  11.38 1.005 12.93 1.235 ;
      RECT  11.38 1.235 11.61 1.565 ;
      RECT  8.23 0.37 9.635 0.6 ;
      RECT  9.405 0.6 9.635 1.565 ;
      RECT  9.14 1.565 11.61 1.795 ;
      RECT  9.965 1.795 10.195 3.53 ;
      RECT  14.95 0.37 15.29 0.6 ;
      RECT  14.95 0.6 15.18 1.005 ;
      RECT  13.83 0.37 14.17 0.6 ;
      RECT  13.94 0.6 14.17 1.005 ;
      RECT  13.16 1.005 15.18 1.235 ;
      RECT  13.16 1.235 13.39 1.565 ;
      RECT  12.765 1.565 13.39 1.795 ;
      RECT  12.765 1.795 12.995 3.245 ;
      RECT  12.765 3.245 13.26 3.475 ;
      RECT  2.42 1.005 5.0 1.235 ;
      RECT  3.96 1.465 8.78 1.695 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 2.405 ;
      RECT  2.685 2.405 4.09 2.635 ;
      RECT  2.685 2.635 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
      RECT  3.245 1.51 3.475 1.925 ;
      RECT  3.245 1.925 7.955 2.155 ;
      RECT  7.725 2.155 7.955 2.405 ;
      RECT  4.365 2.155 4.595 3.03 ;
      RECT  7.725 2.405 9.69 2.635 ;
      RECT  7.725 2.635 7.955 3.245 ;
      RECT  3.19 3.03 4.595 3.26 ;
      RECT  6.9 3.245 7.955 3.475 ;
      RECT  3.96 3.49 5.0 3.72 ;
      RECT  5.46 3.805 10.195 3.95 ;
      RECT  1.565 3.95 10.195 4.035 ;
      RECT  1.565 4.035 5.69 4.18 ;
      RECT  9.965 4.035 10.195 4.925 ;
      RECT  1.565 4.18 1.795 4.365 ;
      RECT  0.18 1.565 0.675 1.795 ;
      RECT  0.445 1.795 0.675 4.365 ;
      RECT  0.18 4.365 1.795 4.595 ;
      RECT  9.965 4.925 11.93 5.155 ;
      RECT  11.59 5.155 11.93 5.23 ;
      RECT  6.045 4.365 8.78 4.41 ;
      RECT  2.42 4.41 8.78 4.595 ;
      RECT  2.42 4.595 6.275 4.64 ;
      RECT  10.68 4.365 11.72 4.595 ;
      RECT  1.51 5.0 2.97 5.23 ;
  END
END MDN_LDPRBSBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_LDPRBSBQ_4
#      Description : D-latch, pos-gate, lo-async-clear, lo-async-set, q-only
#      Equation    : iq,iqn=latch(enable=G,data_in=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDPRBSBQ_4
  CLASS CORE ;
  FOREIGN MDN_LDPRBSBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.915 2.385 5.165 2.66 ;
      RECT  4.925 2.66 5.715 2.94 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.62 1.565 17.74 1.795 ;
      RECT  15.565 1.795 15.795 3.245 ;
      RECT  13.62 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.565 0.37 7.45 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  0.39 0.37 0.73 0.6 ;
      RECT  0.42 0.6 0.7 1.005 ;
      RECT  0.42 1.005 1.795 1.235 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  9.14 4.365 9.635 4.595 ;
      RECT  9.405 4.595 9.635 5.46 ;
      RECT  9.405 5.46 12.435 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  10.525 -0.14 11.2 0.14 ;
      RECT  10.525 0.14 10.755 1.005 ;
      RECT  10.525 1.005 11.02 1.235 ;
      RECT  7.28 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 1.005 ;
      RECT  6.2 1.005 7.955 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.71 0.6 12.94 1.005 ;
      RECT  11.38 1.005 12.94 1.235 ;
      RECT  11.38 1.235 11.61 1.565 ;
      RECT  8.23 0.37 8.57 0.445 ;
      RECT  8.23 0.445 9.33 0.675 ;
      RECT  9.1 0.675 9.33 1.565 ;
      RECT  9.1 1.565 11.61 1.795 ;
      RECT  9.965 1.795 10.195 3.53 ;
      RECT  14.95 0.37 16.41 0.6 ;
      RECT  2.42 1.005 5.0 1.235 ;
      RECT  3.96 1.465 8.78 1.695 ;
      RECT  0.18 1.565 0.675 1.795 ;
      RECT  0.445 1.795 0.675 3.805 ;
      RECT  0.445 3.805 3.475 3.95 ;
      RECT  0.445 3.95 10.195 4.035 ;
      RECT  5.485 3.805 10.195 3.95 ;
      RECT  3.245 4.035 5.715 4.18 ;
      RECT  0.445 4.035 0.675 4.365 ;
      RECT  9.965 4.035 10.195 4.925 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  9.965 4.925 11.93 5.155 ;
      RECT  11.59 5.155 11.93 5.23 ;
      RECT  1.715 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 2.405 ;
      RECT  2.685 2.405 4.09 2.635 ;
      RECT  2.685 2.635 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
      RECT  12.765 1.565 13.26 1.795 ;
      RECT  12.765 1.795 12.995 2.405 ;
      RECT  12.765 2.405 15.29 2.635 ;
      RECT  12.765 2.635 12.995 3.245 ;
      RECT  12.765 3.245 13.26 3.475 ;
      RECT  3.245 1.51 3.475 1.925 ;
      RECT  3.245 1.925 7.955 2.155 ;
      RECT  7.725 2.155 7.955 2.405 ;
      RECT  4.365 2.155 4.595 3.03 ;
      RECT  7.725 2.405 9.69 2.635 ;
      RECT  7.725 2.635 7.955 3.245 ;
      RECT  3.19 3.03 4.595 3.26 ;
      RECT  6.9 3.245 7.955 3.475 ;
      RECT  16.07 2.405 17.53 2.635 ;
      RECT  3.96 3.49 5.0 3.72 ;
      RECT  6.045 4.365 8.78 4.41 ;
      RECT  2.42 4.41 8.78 4.595 ;
      RECT  2.42 4.595 6.275 4.64 ;
      RECT  10.63 4.365 11.72 4.595 ;
      RECT  1.51 5.0 2.97 5.23 ;
  END
END MDN_LDPRBSBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_LDPSBQ_4
#      Description : D-latch, pos-gate, lo-async-set, q-only
#      Equation    : iq,iqn=latch(enable=G,data_in=D,preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDPSBQ_4
  CLASS CORE ;
  FOREIGN MDN_LDPSBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.14 1.565 13.26 1.795 ;
      RECT  11.085 1.795 11.315 3.245 ;
      RECT  9.14 3.245 13.26 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  6.16 -0.14 7.28 0.14 ;
      RECT  6.605 0.14 6.835 1.005 ;
      RECT  6.2 1.005 6.835 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  4.87 0.37 5.21 0.445 ;
      RECT  3.245 0.445 5.21 0.675 ;
      RECT  3.245 0.675 3.475 1.565 ;
      RECT  3.19 1.565 4.43 1.795 ;
      RECT  4.2 1.795 4.43 3.245 ;
      RECT  3.19 3.245 4.43 3.475 ;
      RECT  10.47 0.37 11.93 0.6 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.005 5.715 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  5.485 1.565 7.24 1.795 ;
      RECT  1.72 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 2.405 ;
      RECT  2.125 2.405 3.97 2.635 ;
      RECT  2.125 2.635 2.355 3.245 ;
      RECT  1.72 3.245 2.355 3.475 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 3.245 ;
      RECT  4.66 3.245 6.54 3.475 ;
      RECT  8.285 1.565 8.78 1.795 ;
      RECT  8.285 1.795 8.515 2.405 ;
      RECT  8.285 2.405 10.81 2.635 ;
      RECT  8.285 2.635 8.515 3.245 ;
      RECT  8.285 3.245 8.78 3.475 ;
      RECT  11.59 2.405 13.05 2.635 ;
      RECT  2.42 3.805 7.24 4.035 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  6.2 4.365 8.46 4.595 ;
      RECT  7.22 4.595 7.45 5.0 ;
      RECT  8.23 4.595 8.46 5.0 ;
      RECT  7.11 5.0 7.45 5.23 ;
      RECT  8.23 5.0 8.57 5.23 ;
      RECT  1.51 5.0 2.97 5.23 ;
  END
END MDN_LDPSBQ_4
#-----------------------------------------------------------------------
#      Cell        : MDN_LDPSBQ_1
#      Description : D-latch, pos-gate, lo-async-set, q-only
#      Equation    : iq,iqn=latch(enable=G,data_in=D,preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDPSBQ_1
  CLASS CORE ;
  FOREIGN MDN_LDPSBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.035 2.35 6.285 2.66 ;
      RECT  5.485 2.66 6.275 2.94 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  5.97 0.37 7.45 0.6 ;
      RECT  5.97 0.6 6.2 0.83 ;
      RECT  3.75 0.37 5.23 0.7 ;
      RECT  5.0 0.7 5.23 0.83 ;
      RECT  3.78 0.7 4.06 1.235 ;
      RECT  5.0 0.83 6.2 1.06 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.14 1.005 10.195 1.235 ;
      RECT  9.965 1.235 10.195 4.365 ;
      RECT  9.14 4.365 10.195 4.595 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 2.94 2.355 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  3.19 5.135 3.53 5.46 ;
      RECT  2.8 5.46 6.16 5.74 ;
      RECT  5.43 5.135 5.77 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.6 ;
      RECT  1.68 -0.14 2.8 0.14 ;
      RECT  2.125 0.14 2.355 1.005 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  6.605 1.005 8.78 1.235 ;
      RECT  6.605 1.235 6.835 1.29 ;
      RECT  5.485 1.29 6.835 1.52 ;
      RECT  5.485 1.52 5.715 1.565 ;
      RECT  4.66 1.565 5.715 1.795 ;
      RECT  0.18 1.565 0.52 1.795 ;
      RECT  0.18 1.795 0.41 4.365 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  1.83 4.595 2.06 4.675 ;
      RECT  1.83 4.675 5.09 4.905 ;
      RECT  4.86 4.905 5.09 5.0 ;
      RECT  4.86 5.0 5.2 5.23 ;
      RECT  3.805 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
      RECT  6.2 1.75 7.24 1.98 ;
      RECT  7.725 1.51 7.955 2.685 ;
      RECT  7.725 2.685 9.635 2.915 ;
      RECT  9.405 2.375 9.635 2.685 ;
      RECT  7.725 2.915 7.955 3.705 ;
      RECT  0.64 2.35 0.87 3.705 ;
      RECT  0.64 3.705 7.955 3.935 ;
      RECT  4.66 3.245 7.24 3.475 ;
      RECT  6.2 4.165 6.835 4.365 ;
      RECT  6.2 4.365 8.78 4.395 ;
      RECT  6.605 4.395 8.78 4.595 ;
      RECT  2.42 4.215 5.715 4.445 ;
      RECT  5.485 4.445 5.715 4.63 ;
      RECT  5.485 4.63 6.275 4.86 ;
      RECT  6.045 4.86 6.275 4.925 ;
      RECT  6.045 4.925 8.57 5.155 ;
      RECT  8.23 5.155 8.57 5.23 ;
  END
END MDN_LDPSBQ_1
#-----------------------------------------------------------------------
#      Cell        : MDN_LDPSBQ_2
#      Description : D-latch, pos-gate, lo-async-set, q-only
#      Equation    : iq,iqn=latch(enable=G,data_in=D,preset=!SD):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_LDPSBQ_2
  CLASS CORE ;
  FOREIGN MDN_LDPSBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.63 0.37 5.21 0.6 ;
      RECT  4.9 0.6 5.18 1.235 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.14 1.565 11.025 1.795 ;
      RECT  9.405 1.795 9.635 3.245 ;
      RECT  9.14 3.245 11.02 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 7.42 2.355 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  6.16 -0.14 7.28 0.14 ;
      RECT  6.605 0.14 6.835 1.005 ;
      RECT  6.2 1.005 7.24 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 1.565 ;
      RECT  1.005 1.565 2.76 1.795 ;
      RECT  1.72 1.005 4.3 1.235 ;
      RECT  3.805 1.565 5.0 1.795 ;
      RECT  3.805 1.795 4.035 3.245 ;
      RECT  3.805 3.245 6.54 3.475 ;
      RECT  8.285 1.565 8.78 1.795 ;
      RECT  8.285 1.795 8.515 3.805 ;
      RECT  4.53 3.805 8.78 4.035 ;
      RECT  4.53 4.035 4.76 4.365 ;
      RECT  2.685 4.365 4.76 4.595 ;
      RECT  2.685 4.595 2.915 5.0 ;
      RECT  1.51 5.0 2.915 5.23 ;
      RECT  1.72 3.245 2.76 3.475 ;
      RECT  3.245 1.51 3.475 3.53 ;
      RECT  2.125 3.805 4.3 4.035 ;
      RECT  2.125 4.035 2.355 4.365 ;
      RECT  0.18 4.365 2.355 4.595 ;
      RECT  9.46 4.365 10.7 4.595 ;
      RECT  9.46 4.595 9.69 5.0 ;
      RECT  10.47 4.595 10.7 5.0 ;
      RECT  4.99 4.365 8.46 4.595 ;
      RECT  4.99 4.595 5.22 4.925 ;
      RECT  8.23 4.595 8.46 5.0 ;
      RECT  3.19 4.925 5.22 5.155 ;
      RECT  8.23 5.0 9.69 5.23 ;
      RECT  10.47 5.0 10.81 5.23 ;
  END
END MDN_LDPSBQ_2
#-----------------------------------------------------------------------
#      Cell        : MDN_MAJ3_1
#      Description : 3-input majority
#      Equation    : X=(A1&A2)|(A1&A3)|(A2&A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MAJ3_1
  CLASS CORE ;
  FOREIGN MDN_MAJ3_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 6.89 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 1.565 6.54 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  5.485 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.445 ;
      RECT  1.51 0.445 5.21 0.675 ;
      RECT  4.87 0.37 5.21 0.445 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.245 1.005 6.22 1.235 ;
      RECT  3.245 1.235 3.475 3.53 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.955 1.565 5.0 1.795 ;
      RECT  3.96 3.245 5.0 3.475 ;
      RECT  0.18 3.805 2.76 4.035 ;
      RECT  0.5 4.365 1.795 4.595 ;
      RECT  1.565 4.595 1.795 4.925 ;
      RECT  0.5 4.595 0.73 5.0 ;
      RECT  1.565 4.925 4.09 5.155 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  3.75 5.155 4.09 5.23 ;
  END
END MDN_MAJ3_1
#-----------------------------------------------------------------------
#      Cell        : MDN_MAJ3_2
#      Description : 3-input majority
#      Equation    : X=(A1&A2)|(A1&A3)|(A2&A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MAJ3_2
  CLASS CORE ;
  FOREIGN MDN_MAJ3_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  4.48 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 7.955 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  6.2 3.245 7.955 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.445 ;
      RECT  1.51 0.445 5.21 0.675 ;
      RECT  4.87 0.37 5.21 0.445 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  3.245 1.51 3.475 2.685 ;
      RECT  3.245 2.685 7.395 2.915 ;
      RECT  6.045 2.35 6.275 2.685 ;
      RECT  7.165 2.35 7.395 2.685 ;
      RECT  3.245 2.915 3.475 3.53 ;
      RECT  3.96 3.245 5.0 3.475 ;
      RECT  0.18 3.805 2.355 4.035 ;
      RECT  2.125 4.035 2.355 4.365 ;
      RECT  2.125 4.365 2.76 4.595 ;
      RECT  0.445 4.365 1.795 4.595 ;
      RECT  1.565 4.595 1.795 4.925 ;
      RECT  0.445 4.595 0.675 5.0 ;
      RECT  1.565 4.925 4.09 5.155 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  3.75 5.155 4.09 5.23 ;
  END
END MDN_MAJ3_2
#-----------------------------------------------------------------------
#      Cell        : MDN_MAJ3_4
#      Description : 3-input majority
#      Equation    : X=(A1&A2)|(A1&A3)|(A2&A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MAJ3_4
  CLASS CORE ;
  FOREIGN MDN_MAJ3_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  4.48 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 10.195 1.795 ;
      RECT  9.965 1.795 10.195 3.245 ;
      RECT  6.2 3.245 10.195 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.445 ;
      RECT  1.51 0.445 5.21 0.675 ;
      RECT  4.87 0.37 5.21 0.445 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  3.245 1.585 3.475 2.685 ;
      RECT  3.245 2.685 9.635 2.915 ;
      RECT  6.045 2.35 6.275 2.685 ;
      RECT  7.165 2.35 7.395 2.685 ;
      RECT  8.285 2.35 8.515 2.685 ;
      RECT  9.405 2.35 9.635 2.685 ;
      RECT  3.245 2.915 3.475 3.455 ;
      RECT  3.955 3.245 5.0 3.475 ;
      RECT  0.18 3.805 2.355 4.035 ;
      RECT  2.125 4.035 2.355 4.365 ;
      RECT  2.125 4.365 2.76 4.595 ;
      RECT  0.5 4.365 1.795 4.595 ;
      RECT  1.565 4.595 1.795 4.925 ;
      RECT  0.5 4.595 0.73 5.0 ;
      RECT  1.565 4.925 4.09 5.155 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  3.75 5.155 4.09 5.23 ;
  END
END MDN_MAJ3_4
#-----------------------------------------------------------------------
#      Cell        : MDN_MAJI3_1
#      Description : 3-input majority, inverted
#      Equation    : X=!((A1&A2)|(A1&A3)|(A2&A3))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MAJI3_1
  CLASS CORE ;
  FOREIGN MDN_MAJI3_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 1.51 3.475 3.53 ;
    END
    ANTENNADIFFAREA 2.566 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.445 ;
      RECT  1.51 0.445 5.21 0.675 ;
      RECT  4.87 0.37 5.21 0.445 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  3.96 3.245 5.0 3.475 ;
      RECT  0.18 3.805 2.76 4.035 ;
      RECT  0.5 4.365 1.795 4.595 ;
      RECT  1.565 4.595 1.795 4.925 ;
      RECT  0.5 4.595 0.73 5.0 ;
      RECT  1.565 4.925 4.09 5.155 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  3.75 5.155 4.09 5.23 ;
  END
END MDN_MAJI3_1
#-----------------------------------------------------------------------
#      Cell        : MDN_MAJI3_2
#      Description : 3-input majority, inverted
#      Equation    : X=!((A1&A2)|(A1&A3)|(A2&A3))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MAJI3_2
  CLASS CORE ;
  FOREIGN MDN_MAJI3_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 10.78 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 5.46 11.37 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 -0.14 11.37 0.14 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.895 1.005 11.02 1.235 ;
      RECT  8.845 1.235 9.075 4.365 ;
      RECT  6.895 4.365 11.02 4.595 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  6.31 0.445 10.25 0.675 ;
      RECT  6.31 0.675 6.54 1.005 ;
      RECT  2.42 1.005 6.54 1.235 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 8.01 1.795 ;
      RECT  1.565 3.805 8.01 4.035 ;
      RECT  1.565 4.035 1.795 4.365 ;
      RECT  0.18 4.365 1.795 4.595 ;
      RECT  2.42 4.365 6.54 4.595 ;
      RECT  6.31 4.595 6.54 4.925 ;
      RECT  6.31 4.925 10.25 5.155 ;
  END
END MDN_MAJI3_2
#-----------------------------------------------------------------------
#      Cell        : MDN_MAJI3_4
#      Description : 3-input majority, inverted
#      Equation    : X=!((A1&A2)|(A1&A3)|(A2&A3))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MAJI3_4
  CLASS CORE ;
  FOREIGN MDN_MAJI3_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 17.5 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 4.536 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 8.54 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 4.536 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.34 2.125 21.98 2.355 ;
      RECT  18.34 2.355 18.62 2.915 ;
      RECT  19.46 2.355 19.74 2.915 ;
      RECT  20.58 2.355 20.86 2.915 ;
      RECT  21.7 2.355 21.98 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.84 5.46 22.57 5.74 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.84 -0.14 22.57 0.14 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.62 1.005 22.22 1.235 ;
      RECT  17.805 1.235 18.035 4.365 ;
      RECT  13.62 4.365 22.22 4.595 ;
    END
    ANTENNADIFFAREA 12.096 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  13.03 0.445 21.45 0.675 ;
      RECT  13.03 0.675 13.26 1.005 ;
      RECT  4.66 1.005 13.26 1.235 ;
      RECT  0.18 1.005 4.035 1.235 ;
      RECT  3.805 1.235 4.035 1.565 ;
      RECT  3.805 1.565 16.97 1.795 ;
      RECT  3.805 3.805 16.97 4.035 ;
      RECT  3.805 4.035 4.035 4.365 ;
      RECT  0.18 4.365 4.035 4.595 ;
      RECT  4.66 4.365 13.26 4.595 ;
      RECT  13.03 4.595 13.26 4.925 ;
      RECT  13.03 4.925 21.45 5.155 ;
  END
END MDN_MAJI3_4
#-----------------------------------------------------------------------
#      Cell        : MDN_MUX2_1
#      Description : 2-1 multiplexer
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUX2_1
  CLASS CORE ;
  FOREIGN MDN_MUX2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  6.16 5.46 6.89 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  4.31 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  1.005 5.46 1.68 5.74 ;
      RECT  -0.17 5.46 0.56 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  6.16 -0.14 6.89 0.14 ;
      RECT  4.31 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  1.565 -0.14 2.41 0.14 ;
      RECT  1.565 0.14 1.795 1.005 ;
      RECT  1.565 1.005 2.76 1.235 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.245 1.005 6.22 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 1.565 ;
      RECT  1.005 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 3.53 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 4.365 ;
      RECT  4.66 4.365 5.155 4.595 ;
      RECT  4.925 4.595 5.155 4.925 ;
      RECT  1.51 4.925 5.155 5.155 ;
      RECT  1.51 5.155 1.85 5.23 ;
      RECT  0.18 4.365 4.3 4.595 ;
  END
END MDN_MUX2_1
#-----------------------------------------------------------------------
#      Cell        : MDN_MUX2_2
#      Description : 2-1 multiplexer
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUX2_2
  CLASS CORE ;
  FOREIGN MDN_MUX2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 9.13 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  4.31 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  8.4 -0.14 9.13 0.14 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  4.31 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  1.68 -0.14 2.8 0.14 ;
      RECT  2.125 0.14 2.355 1.005 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  6.2 3.245 7.24 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.245 1.005 6.22 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 1.565 ;
      RECT  1.005 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 3.53 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 4.365 ;
      RECT  4.66 4.365 5.155 4.595 ;
      RECT  4.925 4.595 5.155 4.925 ;
      RECT  1.51 4.925 5.155 5.155 ;
      RECT  1.51 5.155 1.85 5.23 ;
      RECT  0.18 4.365 4.3 4.595 ;
  END
END MDN_MUX2_2
#-----------------------------------------------------------------------
#      Cell        : MDN_MUX2_3
#      Description : 2-1 multiplexer
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUX2_3
  CLASS CORE ;
  FOREIGN MDN_MUX2_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 9.13 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  4.31 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  8.4 -0.14 9.13 0.14 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  1.565 -0.14 2.41 0.14 ;
      RECT  1.565 0.14 1.795 1.005 ;
      RECT  1.565 1.005 2.76 1.235 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 8.78 1.795 ;
      RECT  7.165 1.795 7.395 3.245 ;
      RECT  6.2 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 4.536 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  8.23 0.37 8.57 0.6 ;
      RECT  8.23 0.6 8.46 1.005 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  7.22 0.6 7.45 1.005 ;
      RECT  3.245 1.005 6.22 1.235 ;
      RECT  7.22 1.005 8.46 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 1.565 ;
      RECT  1.005 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 3.53 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 4.365 ;
      RECT  4.66 4.365 5.155 4.595 ;
      RECT  4.925 4.595 5.155 4.925 ;
      RECT  1.51 4.925 5.155 5.155 ;
      RECT  1.51 5.155 1.85 5.23 ;
      RECT  0.18 4.365 4.3 4.595 ;
  END
END MDN_MUX2_3
#-----------------------------------------------------------------------
#      Cell        : MDN_MUX2_4
#      Description : 2-1 multiplexer
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUX2_4
  CLASS CORE ;
  FOREIGN MDN_MUX2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.905 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.905 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.905 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.905 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  1.68 -0.14 2.8 0.14 ;
      RECT  2.125 0.14 2.355 1.005 ;
      RECT  1.72 1.005 2.76 1.235 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 9.48 1.795 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  6.2 3.245 9.48 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  8.23 0.37 9.69 0.6 ;
      RECT  3.245 1.005 5.715 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  5.485 1.235 5.715 2.405 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 1.565 ;
      RECT  1.005 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 3.455 ;
      RECT  5.485 2.405 8.57 2.635 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 4.365 ;
      RECT  4.66 4.365 5.155 4.595 ;
      RECT  4.925 4.595 5.155 5.0 ;
      RECT  1.51 5.0 5.155 5.23 ;
      RECT  0.18 4.365 4.3 4.595 ;
  END
END MDN_MUX2_4
#-----------------------------------------------------------------------
#      Cell        : MDN_MUX2B_1
#      Description : 2-1 multiplexer with D0 input inverted
#      Equation    : X=(S&D1)|(!S&!D0)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUX2B_1
  CLASS CORE ;
  FOREIGN MDN_MUX2B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 4.365 1.795 4.595 ;
      RECT  0.42 4.595 0.7 5.0 ;
      RECT  1.565 4.595 1.795 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  1.565 5.0 6.33 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.43 4.365 6.835 4.595 ;
      RECT  6.605 4.595 6.835 5.46 ;
      RECT  6.16 5.46 7.955 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 7.955 1.795 ;
      RECT  7.725 1.795 7.955 3.805 ;
      RECT  6.9 3.805 7.955 4.035 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.565 0.37 5.21 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  0.445 1.235 0.675 3.245 ;
      RECT  0.18 3.245 0.675 3.475 ;
      RECT  2.42 1.005 5.0 1.235 ;
      RECT  5.49 1.005 6.54 1.235 ;
      RECT  5.49 1.235 5.72 1.565 ;
      RECT  3.96 1.565 5.72 1.795 ;
      RECT  1.7 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.805 ;
      RECT  1.72 3.805 2.915 4.035 ;
      RECT  3.245 1.51 3.475 3.245 ;
      RECT  3.245 3.245 7.395 3.475 ;
      RECT  7.165 2.35 7.395 3.245 ;
      RECT  3.245 3.805 6.54 4.035 ;
      RECT  3.245 4.035 3.475 4.365 ;
      RECT  2.42 4.365 3.475 4.595 ;
      RECT  3.96 4.365 5.0 4.595 ;
  END
END MDN_MUX2B_1
#-----------------------------------------------------------------------
#      Cell        : MDN_MUX2B_2
#      Description : 2-1 multiplexer with D0 input inverted
#      Equation    : X=(S&D1)|(!S&!D0)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUX2B_2
  CLASS CORE ;
  FOREIGN MDN_MUX2B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 4.365 1.795 4.595 ;
      RECT  0.42 4.595 0.7 5.0 ;
      RECT  1.565 4.595 1.795 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  1.565 5.0 6.33 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.43 4.365 6.835 4.595 ;
      RECT  6.605 4.595 6.835 5.46 ;
      RECT  6.16 5.46 7.955 5.74 ;
      RECT  7.725 4.905 7.955 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 8.78 1.795 ;
      RECT  7.725 1.795 7.955 3.805 ;
      RECT  6.9 3.805 8.78 4.035 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.565 0.37 5.21 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  0.445 1.235 0.675 3.245 ;
      RECT  0.18 3.245 0.675 3.475 ;
      RECT  2.42 1.005 5.0 1.235 ;
      RECT  5.49 1.005 6.54 1.235 ;
      RECT  5.49 1.235 5.72 1.565 ;
      RECT  3.96 1.565 5.72 1.795 ;
      RECT  1.7 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.805 ;
      RECT  1.72 3.805 2.915 4.035 ;
      RECT  3.245 1.51 3.475 3.245 ;
      RECT  3.245 3.245 7.395 3.475 ;
      RECT  7.165 2.35 7.395 3.245 ;
      RECT  3.245 3.805 6.54 4.035 ;
      RECT  3.245 4.035 3.475 4.365 ;
      RECT  2.42 4.365 3.475 4.595 ;
      RECT  3.96 4.365 5.0 4.595 ;
      RECT  7.22 4.365 8.46 4.595 ;
      RECT  7.22 4.595 7.45 5.0 ;
      RECT  8.23 4.595 8.46 5.0 ;
      RECT  7.11 5.0 7.45 5.23 ;
      RECT  8.23 5.0 8.57 5.23 ;
  END
END MDN_MUX2B_2
#-----------------------------------------------------------------------
#      Cell        : MDN_MUX2B_3
#      Description : 2-1 multiplexer with D0 input inverted
#      Equation    : X=(S&D1)|(!S&!D0)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUX2B_3
  CLASS CORE ;
  FOREIGN MDN_MUX2B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 4.365 1.795 4.595 ;
      RECT  0.42 4.595 0.7 5.0 ;
      RECT  1.565 4.595 1.795 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  1.565 5.0 6.33 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.905 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  5.43 4.365 6.835 4.595 ;
      RECT  6.605 4.595 6.835 5.46 ;
      RECT  6.16 5.46 7.955 5.74 ;
      RECT  7.725 4.905 7.955 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 9.48 1.795 ;
      RECT  8.845 1.795 9.075 3.805 ;
      RECT  6.9 3.805 9.48 4.035 ;
    END
    ANTENNADIFFAREA 4.536 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.565 0.37 5.21 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  0.445 1.235 0.675 3.245 ;
      RECT  0.18 3.245 0.675 3.475 ;
      RECT  2.42 1.005 5.0 1.235 ;
      RECT  5.49 1.005 6.54 1.235 ;
      RECT  5.49 1.235 5.72 1.565 ;
      RECT  3.96 1.565 5.72 1.795 ;
      RECT  1.7 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.805 ;
      RECT  1.72 3.805 2.915 4.035 ;
      RECT  7.165 2.405 8.43 2.635 ;
      RECT  7.165 2.635 7.395 3.245 ;
      RECT  3.245 1.51 3.475 3.245 ;
      RECT  3.245 3.245 7.395 3.475 ;
      RECT  3.245 3.805 6.54 4.035 ;
      RECT  3.245 4.035 3.475 4.365 ;
      RECT  2.42 4.365 3.475 4.595 ;
      RECT  3.96 4.365 5.0 4.595 ;
      RECT  8.23 5.0 9.69 5.23 ;
  END
END MDN_MUX2B_3
#-----------------------------------------------------------------------
#      Cell        : MDN_MUX2B_4
#      Description : 2-1 multiplexer with D0 input inverted
#      Equation    : X=(S&D1)|(!S&!D0)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUX2B_4
  CLASS CORE ;
  FOREIGN MDN_MUX2B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 4.365 1.795 4.595 ;
      RECT  0.42 4.595 0.7 5.0 ;
      RECT  1.565 4.595 1.795 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
      RECT  1.565 5.0 6.33 5.23 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.905 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  5.43 4.365 6.835 4.595 ;
      RECT  6.605 4.595 6.835 5.46 ;
      RECT  6.16 5.46 7.955 5.74 ;
      RECT  7.725 4.905 7.955 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 11.02 1.795 ;
      RECT  9.965 1.795 10.195 3.805 ;
      RECT  6.9 3.805 11.02 4.035 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.565 0.37 5.21 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  0.445 1.235 0.675 3.245 ;
      RECT  0.18 3.245 0.675 3.475 ;
      RECT  2.42 1.005 5.0 1.235 ;
      RECT  5.49 1.005 6.54 1.235 ;
      RECT  5.49 1.235 5.72 1.565 ;
      RECT  3.96 1.565 5.72 1.795 ;
      RECT  1.7 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.805 ;
      RECT  1.72 3.805 2.915 4.035 ;
      RECT  7.165 2.405 9.545 2.635 ;
      RECT  7.165 2.635 7.395 3.245 ;
      RECT  3.245 1.51 3.475 3.245 ;
      RECT  3.245 3.245 7.395 3.475 ;
      RECT  3.245 3.805 6.54 4.035 ;
      RECT  3.245 4.035 3.475 4.365 ;
      RECT  2.42 4.365 3.475 4.595 ;
      RECT  3.96 4.365 5.0 4.595 ;
      RECT  9.46 4.365 10.7 4.595 ;
      RECT  9.46 4.595 9.69 5.0 ;
      RECT  10.47 4.595 10.7 5.0 ;
      RECT  9.35 5.0 9.69 5.23 ;
      RECT  10.47 5.0 10.81 5.23 ;
  END
END MDN_MUX2B_4
#-----------------------------------------------------------------------
#      Cell        : MDN_MUX4_1
#      Description : 4-1 multiplexer
#      Equation    : X=((D0&!S0&!S1)|(D1&S0&!S1)|(D2&!S0&S1)|(D3&S0&S1))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUX4_1
  CLASS CORE ;
  FOREIGN MDN_MUX4_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D2
  PIN D3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D3
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 14.14 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.87 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 10.64 5.74 ;
      RECT  3.245 5.065 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  9.52 -0.14 10.64 0.14 ;
      RECT  9.91 0.14 10.25 0.465 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 1.005 ;
      RECT  1.005 1.005 3.53 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 3.245 ;
      RECT  15.005 3.245 15.5 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.445 ;
      RECT  1.51 0.445 7.45 0.675 ;
      RECT  4.87 0.37 5.21 0.445 ;
      RECT  7.11 0.37 7.45 0.445 ;
      RECT  11.59 0.37 14.17 0.6 ;
      RECT  7.725 0.695 10.195 0.925 ;
      RECT  7.725 0.925 7.955 1.005 ;
      RECT  9.965 0.925 10.195 1.005 ;
      RECT  6.9 1.005 7.955 1.235 ;
      RECT  9.965 1.005 11.02 1.235 ;
      RECT  12.21 1.005 13.26 1.01 ;
      RECT  12.205 1.01 13.26 1.015 ;
      RECT  12.2 1.015 13.26 1.02 ;
      RECT  12.195 1.02 13.26 1.025 ;
      RECT  12.19 1.025 13.26 1.03 ;
      RECT  12.185 1.03 13.26 1.035 ;
      RECT  12.18 1.035 13.26 1.04 ;
      RECT  12.175 1.04 13.26 1.045 ;
      RECT  12.17 1.045 13.26 1.05 ;
      RECT  12.165 1.05 13.26 1.055 ;
      RECT  12.16 1.055 13.26 1.06 ;
      RECT  12.155 1.06 13.26 1.065 ;
      RECT  12.15 1.065 13.26 1.07 ;
      RECT  12.145 1.07 13.26 1.075 ;
      RECT  12.14 1.075 13.26 1.08 ;
      RECT  12.135 1.08 13.26 1.085 ;
      RECT  12.13 1.085 13.26 1.09 ;
      RECT  12.125 1.09 13.26 1.095 ;
      RECT  12.12 1.095 13.26 1.1 ;
      RECT  12.115 1.1 13.26 1.105 ;
      RECT  12.11 1.105 13.26 1.11 ;
      RECT  12.105 1.11 13.26 1.115 ;
      RECT  12.1 1.115 13.26 1.12 ;
      RECT  12.095 1.12 13.26 1.125 ;
      RECT  12.09 1.125 13.26 1.13 ;
      RECT  12.085 1.13 13.26 1.135 ;
      RECT  12.08 1.135 13.26 1.14 ;
      RECT  12.075 1.14 13.26 1.145 ;
      RECT  12.07 1.145 13.26 1.15 ;
      RECT  12.065 1.15 13.26 1.155 ;
      RECT  12.06 1.155 13.26 1.16 ;
      RECT  12.055 1.16 13.26 1.165 ;
      RECT  12.05 1.165 13.26 1.17 ;
      RECT  12.045 1.17 13.26 1.175 ;
      RECT  12.04 1.175 13.26 1.18 ;
      RECT  12.035 1.18 13.26 1.185 ;
      RECT  12.03 1.185 13.26 1.19 ;
      RECT  12.025 1.19 13.26 1.195 ;
      RECT  12.02 1.195 13.26 1.2 ;
      RECT  12.015 1.2 13.26 1.205 ;
      RECT  12.01 1.205 13.26 1.21 ;
      RECT  12.005 1.21 13.26 1.215 ;
      RECT  12.0 1.215 13.26 1.22 ;
      RECT  11.995 1.22 13.26 1.225 ;
      RECT  11.99 1.225 13.26 1.23 ;
      RECT  11.985 1.23 13.26 1.235 ;
      RECT  11.98 1.235 12.305 1.24 ;
      RECT  11.975 1.24 12.3 1.245 ;
      RECT  11.97 1.245 12.295 1.25 ;
      RECT  11.965 1.25 12.29 1.255 ;
      RECT  11.96 1.255 12.285 1.26 ;
      RECT  11.955 1.26 12.28 1.265 ;
      RECT  11.95 1.265 12.275 1.27 ;
      RECT  11.945 1.27 12.27 1.275 ;
      RECT  11.94 1.275 12.265 1.28 ;
      RECT  11.935 1.28 12.26 1.285 ;
      RECT  11.93 1.285 12.255 1.29 ;
      RECT  11.925 1.29 12.25 1.295 ;
      RECT  11.92 1.295 12.245 1.3 ;
      RECT  11.915 1.3 12.24 1.305 ;
      RECT  11.91 1.305 12.235 1.31 ;
      RECT  11.905 1.31 12.23 1.315 ;
      RECT  11.9 1.315 12.225 1.32 ;
      RECT  11.895 1.32 12.22 1.325 ;
      RECT  11.89 1.325 12.215 1.33 ;
      RECT  11.885 1.33 12.21 1.335 ;
      RECT  11.88 1.335 12.205 1.34 ;
      RECT  11.875 1.34 12.2 1.345 ;
      RECT  11.87 1.345 12.195 1.35 ;
      RECT  11.865 1.35 12.19 1.355 ;
      RECT  11.86 1.355 12.185 1.36 ;
      RECT  11.855 1.36 12.18 1.365 ;
      RECT  11.85 1.365 12.175 1.37 ;
      RECT  11.845 1.37 12.17 1.375 ;
      RECT  11.84 1.375 12.165 1.38 ;
      RECT  11.835 1.38 12.16 1.385 ;
      RECT  11.83 1.385 12.155 1.39 ;
      RECT  11.825 1.39 12.15 1.395 ;
      RECT  11.82 1.395 12.145 1.4 ;
      RECT  11.815 1.4 12.14 1.405 ;
      RECT  11.81 1.405 12.135 1.41 ;
      RECT  11.805 1.41 12.13 1.415 ;
      RECT  11.8 1.415 12.125 1.42 ;
      RECT  11.795 1.42 12.12 1.425 ;
      RECT  11.79 1.425 12.115 1.43 ;
      RECT  11.785 1.43 12.11 1.435 ;
      RECT  11.78 1.435 12.105 1.44 ;
      RECT  11.775 1.44 12.1 1.445 ;
      RECT  11.77 1.445 12.095 1.45 ;
      RECT  11.765 1.45 12.09 1.455 ;
      RECT  11.76 1.455 12.085 1.46 ;
      RECT  11.755 1.46 12.08 1.465 ;
      RECT  11.75 1.465 12.075 1.47 ;
      RECT  11.745 1.47 12.07 1.475 ;
      RECT  11.745 1.475 12.065 1.48 ;
      RECT  11.745 1.48 12.06 1.485 ;
      RECT  11.745 1.485 12.055 1.49 ;
      RECT  11.745 1.49 12.05 1.495 ;
      RECT  11.745 1.495 12.045 1.5 ;
      RECT  11.745 1.5 12.04 1.505 ;
      RECT  11.745 1.505 12.035 1.51 ;
      RECT  11.745 1.51 12.03 1.515 ;
      RECT  11.745 1.515 12.025 1.52 ;
      RECT  11.745 1.52 12.02 1.525 ;
      RECT  11.745 1.525 12.015 1.53 ;
      RECT  11.745 1.53 12.01 1.535 ;
      RECT  11.745 1.535 12.005 1.54 ;
      RECT  11.745 1.54 12.0 1.545 ;
      RECT  11.745 1.545 11.995 1.55 ;
      RECT  11.745 1.55 11.99 1.555 ;
      RECT  11.745 1.555 11.985 1.56 ;
      RECT  11.745 1.56 11.98 1.565 ;
      RECT  11.745 1.565 11.975 3.245 ;
      RECT  11.38 3.245 11.975 3.475 ;
      RECT  11.275 0.89 11.72 1.12 ;
      RECT  11.275 1.12 11.505 1.565 ;
      RECT  9.965 1.565 11.505 1.615 ;
      RECT  7.67 1.615 11.505 1.795 ;
      RECT  7.67 1.795 10.195 1.845 ;
      RECT  8.845 1.845 9.075 3.245 ;
      RECT  7.67 3.245 10.195 3.475 ;
      RECT  9.965 3.475 10.195 3.705 ;
      RECT  9.965 3.705 12.435 3.935 ;
      RECT  12.205 3.935 12.435 4.365 ;
      RECT  12.205 4.365 13.26 4.595 ;
      RECT  3.96 1.005 6.54 1.235 ;
      RECT  8.44 1.155 9.48 1.385 ;
      RECT  0.18 1.565 1.235 1.795 ;
      RECT  1.005 1.795 1.235 4.365 ;
      RECT  0.18 4.365 1.74 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 2.245 4.035 ;
      RECT  2.015 4.035 2.245 4.605 ;
      RECT  2.015 4.605 4.035 4.835 ;
      RECT  3.805 4.835 4.035 5.0 ;
      RECT  3.805 5.0 6.33 5.23 ;
      RECT  2.42 1.565 5.0 1.795 ;
      RECT  13.325 1.565 13.96 1.795 ;
      RECT  13.325 1.795 13.555 2.405 ;
      RECT  12.71 2.405 13.555 2.635 ;
      RECT  13.325 2.635 13.555 3.245 ;
      RECT  13.325 3.245 13.96 3.475 ;
      RECT  5.99 2.405 8.57 2.635 ;
      RECT  12.205 1.695 12.435 3.245 ;
      RECT  12.205 3.245 12.995 3.475 ;
      RECT  12.765 3.475 12.995 3.805 ;
      RECT  12.765 3.805 14.115 4.035 ;
      RECT  13.885 4.035 14.115 4.365 ;
      RECT  13.885 4.365 15.18 4.595 ;
      RECT  14.95 4.595 15.18 5.0 ;
      RECT  14.95 5.0 15.29 5.23 ;
      RECT  5.485 1.51 5.715 3.455 ;
      RECT  2.475 3.685 6.54 3.915 ;
      RECT  2.475 3.915 2.705 4.09 ;
      RECT  6.9 3.705 9.48 3.935 ;
      RECT  3.96 4.145 5.0 4.375 ;
      RECT  8.44 4.165 11.02 4.395 ;
      RECT  5.43 4.365 7.955 4.595 ;
      RECT  7.725 4.595 7.955 4.625 ;
      RECT  7.725 4.625 11.665 4.855 ;
      RECT  11.435 4.425 11.665 4.625 ;
  END
END MDN_MUX4_1
#-----------------------------------------------------------------------
#      Cell        : MDN_MUX4_2
#      Description : 4-1 multiplexer
#      Equation    : X=((D0&!S0&!S1)|(D1&S0&!S1)|(D2&!S0&S1)|(D3&S0&S1))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUX4_2
  CLASS CORE ;
  FOREIGN MDN_MUX4_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D2
  PIN D3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D3
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 14.14 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.93 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.93 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 10.64 5.74 ;
      RECT  3.245 4.905 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  9.52 -0.14 10.64 0.14 ;
      RECT  9.91 0.14 10.25 0.465 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 1.005 ;
      RECT  1.005 1.005 3.53 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.16 1.565 16.2 1.795 ;
      RECT  15.565 1.795 15.795 3.245 ;
      RECT  15.16 3.245 16.2 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.445 ;
      RECT  1.51 0.445 7.45 0.675 ;
      RECT  4.87 0.37 5.21 0.445 ;
      RECT  7.11 0.37 7.45 0.445 ;
      RECT  11.59 0.37 14.17 0.6 ;
      RECT  7.725 0.695 10.195 0.905 ;
      RECT  6.9 0.905 10.195 0.925 ;
      RECT  9.965 0.925 10.195 1.005 ;
      RECT  6.9 0.925 7.955 1.135 ;
      RECT  9.965 1.005 11.02 1.235 ;
      RECT  12.22 1.005 13.26 1.01 ;
      RECT  12.215 1.01 13.26 1.015 ;
      RECT  12.21 1.015 13.26 1.02 ;
      RECT  12.205 1.02 13.26 1.025 ;
      RECT  12.2 1.025 13.26 1.03 ;
      RECT  12.195 1.03 13.26 1.035 ;
      RECT  12.19 1.035 13.26 1.04 ;
      RECT  12.185 1.04 13.26 1.045 ;
      RECT  12.18 1.045 13.26 1.05 ;
      RECT  12.175 1.05 13.26 1.055 ;
      RECT  12.17 1.055 13.26 1.06 ;
      RECT  12.165 1.06 13.26 1.065 ;
      RECT  12.16 1.065 13.26 1.07 ;
      RECT  12.155 1.07 13.26 1.075 ;
      RECT  12.15 1.075 13.26 1.08 ;
      RECT  12.145 1.08 13.26 1.085 ;
      RECT  12.14 1.085 13.26 1.09 ;
      RECT  12.135 1.09 13.26 1.095 ;
      RECT  12.13 1.095 13.26 1.1 ;
      RECT  12.125 1.1 13.26 1.105 ;
      RECT  12.12 1.105 13.26 1.11 ;
      RECT  12.115 1.11 13.26 1.115 ;
      RECT  12.11 1.115 13.26 1.12 ;
      RECT  12.105 1.12 13.26 1.125 ;
      RECT  12.1 1.125 13.26 1.13 ;
      RECT  12.095 1.13 13.26 1.135 ;
      RECT  12.09 1.135 13.26 1.14 ;
      RECT  12.085 1.14 13.26 1.145 ;
      RECT  12.08 1.145 13.26 1.15 ;
      RECT  12.075 1.15 13.26 1.155 ;
      RECT  12.07 1.155 13.26 1.16 ;
      RECT  12.065 1.16 13.26 1.165 ;
      RECT  12.06 1.165 13.26 1.17 ;
      RECT  12.055 1.17 13.26 1.175 ;
      RECT  12.05 1.175 13.26 1.18 ;
      RECT  12.045 1.18 13.26 1.185 ;
      RECT  12.04 1.185 13.26 1.19 ;
      RECT  12.035 1.19 13.26 1.195 ;
      RECT  12.03 1.195 13.26 1.2 ;
      RECT  12.025 1.2 13.26 1.205 ;
      RECT  12.02 1.205 13.26 1.21 ;
      RECT  12.015 1.21 13.26 1.215 ;
      RECT  12.01 1.215 13.26 1.22 ;
      RECT  12.005 1.22 13.26 1.225 ;
      RECT  12.0 1.225 13.26 1.23 ;
      RECT  11.995 1.23 13.26 1.235 ;
      RECT  11.99 1.235 12.315 1.24 ;
      RECT  11.985 1.24 12.31 1.245 ;
      RECT  11.98 1.245 12.305 1.25 ;
      RECT  11.975 1.25 12.3 1.255 ;
      RECT  11.97 1.255 12.295 1.26 ;
      RECT  11.965 1.26 12.29 1.265 ;
      RECT  11.96 1.265 12.285 1.27 ;
      RECT  11.955 1.27 12.28 1.275 ;
      RECT  11.95 1.275 12.275 1.28 ;
      RECT  11.945 1.28 12.27 1.285 ;
      RECT  11.94 1.285 12.265 1.29 ;
      RECT  11.935 1.29 12.26 1.295 ;
      RECT  11.93 1.295 12.255 1.3 ;
      RECT  11.925 1.3 12.25 1.305 ;
      RECT  11.92 1.305 12.245 1.31 ;
      RECT  11.915 1.31 12.24 1.315 ;
      RECT  11.91 1.315 12.235 1.32 ;
      RECT  11.905 1.32 12.23 1.325 ;
      RECT  11.9 1.325 12.225 1.33 ;
      RECT  11.895 1.33 12.22 1.335 ;
      RECT  11.89 1.335 12.215 1.34 ;
      RECT  11.885 1.34 12.21 1.345 ;
      RECT  11.88 1.345 12.205 1.35 ;
      RECT  11.875 1.35 12.2 1.355 ;
      RECT  11.87 1.355 12.195 1.36 ;
      RECT  11.865 1.36 12.19 1.365 ;
      RECT  11.86 1.365 12.185 1.37 ;
      RECT  11.855 1.37 12.18 1.375 ;
      RECT  11.85 1.375 12.175 1.38 ;
      RECT  11.845 1.38 12.17 1.385 ;
      RECT  11.84 1.385 12.165 1.39 ;
      RECT  11.835 1.39 12.16 1.395 ;
      RECT  11.83 1.395 12.155 1.4 ;
      RECT  11.825 1.4 12.15 1.405 ;
      RECT  11.82 1.405 12.145 1.41 ;
      RECT  11.815 1.41 12.14 1.415 ;
      RECT  11.81 1.415 12.135 1.42 ;
      RECT  11.805 1.42 12.13 1.425 ;
      RECT  11.8 1.425 12.125 1.43 ;
      RECT  11.795 1.43 12.12 1.435 ;
      RECT  11.79 1.435 12.115 1.44 ;
      RECT  11.785 1.44 12.11 1.445 ;
      RECT  11.78 1.445 12.105 1.45 ;
      RECT  11.775 1.45 12.1 1.455 ;
      RECT  11.77 1.455 12.095 1.46 ;
      RECT  11.765 1.46 12.09 1.465 ;
      RECT  11.76 1.465 12.085 1.47 ;
      RECT  11.755 1.47 12.08 1.475 ;
      RECT  11.75 1.475 12.075 1.48 ;
      RECT  11.745 1.48 12.07 1.485 ;
      RECT  11.74 1.485 12.065 1.49 ;
      RECT  11.735 1.49 12.06 1.495 ;
      RECT  11.735 1.495 12.055 1.5 ;
      RECT  11.735 1.5 12.05 1.505 ;
      RECT  11.735 1.505 12.045 1.51 ;
      RECT  11.735 1.51 12.04 1.515 ;
      RECT  11.735 1.515 12.035 1.52 ;
      RECT  11.735 1.52 12.03 1.525 ;
      RECT  11.735 1.525 12.025 1.53 ;
      RECT  11.735 1.53 12.02 1.535 ;
      RECT  11.735 1.535 12.015 1.54 ;
      RECT  11.735 1.54 12.01 1.545 ;
      RECT  11.735 1.545 12.005 1.55 ;
      RECT  11.735 1.55 12.0 1.555 ;
      RECT  11.735 1.555 11.995 1.56 ;
      RECT  11.735 1.56 11.99 1.565 ;
      RECT  11.735 1.565 11.985 1.57 ;
      RECT  11.735 1.57 11.98 1.575 ;
      RECT  11.735 1.575 11.975 1.58 ;
      RECT  11.735 1.58 11.97 1.585 ;
      RECT  11.735 1.585 11.965 3.245 ;
      RECT  11.38 3.245 11.965 3.475 ;
      RECT  11.275 0.89 11.72 1.12 ;
      RECT  11.275 1.12 11.505 1.615 ;
      RECT  7.67 1.615 11.505 1.845 ;
      RECT  8.845 1.845 9.075 3.245 ;
      RECT  7.67 3.245 10.195 3.475 ;
      RECT  9.965 3.475 10.195 3.755 ;
      RECT  9.965 3.755 12.41 3.985 ;
      RECT  12.18 3.985 12.41 4.365 ;
      RECT  12.18 4.365 13.26 4.595 ;
      RECT  3.96 1.005 6.54 1.235 ;
      RECT  8.44 1.155 9.48 1.385 ;
      RECT  0.18 1.565 1.235 1.795 ;
      RECT  1.005 1.795 1.235 4.365 ;
      RECT  0.18 4.365 1.74 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 2.245 4.035 ;
      RECT  2.015 4.035 2.245 4.365 ;
      RECT  2.015 4.365 4.035 4.595 ;
      RECT  3.805 4.595 4.035 5.0 ;
      RECT  3.805 5.0 6.33 5.23 ;
      RECT  2.42 1.565 5.0 1.795 ;
      RECT  13.325 1.565 13.96 1.795 ;
      RECT  13.325 1.795 13.555 2.405 ;
      RECT  12.71 2.405 13.555 2.635 ;
      RECT  13.325 2.635 13.555 3.245 ;
      RECT  13.325 3.245 13.96 3.475 ;
      RECT  5.99 2.405 8.57 2.635 ;
      RECT  12.205 1.695 12.435 3.245 ;
      RECT  12.205 3.245 12.995 3.475 ;
      RECT  12.765 3.475 12.995 3.805 ;
      RECT  12.765 3.805 14.115 4.035 ;
      RECT  13.885 4.035 14.115 4.365 ;
      RECT  13.885 4.365 15.18 4.595 ;
      RECT  14.95 4.595 15.18 5.0 ;
      RECT  14.95 5.0 16.41 5.23 ;
      RECT  5.485 1.51 5.715 3.455 ;
      RECT  3.96 3.245 5.0 3.475 ;
      RECT  6.9 3.705 9.48 3.935 ;
      RECT  6.9 3.935 7.24 4.03 ;
      RECT  2.475 3.795 6.54 4.025 ;
      RECT  2.475 4.025 2.705 4.135 ;
      RECT  8.44 4.215 11.02 4.445 ;
      RECT  5.43 4.365 7.955 4.595 ;
      RECT  7.725 4.595 7.955 4.675 ;
      RECT  7.725 4.675 11.72 4.905 ;
      RECT  11.38 4.48 11.72 4.675 ;
  END
END MDN_MUX4_2
#-----------------------------------------------------------------------
#      Cell        : MDN_MUX4_4
#      Description : 4-1 multiplexer
#      Equation    : X=((D0&!S0&!S1)|(D1&S0&!S1)|(D2&!S0&S1)|(D3&S0&S1))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUX4_4
  CLASS CORE ;
  FOREIGN MDN_MUX4_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D2
  PIN D3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D3
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 14.14 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.93 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  14.445 4.87 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 11.76 5.74 ;
      RECT  3.245 5.08 3.475 5.46 ;
      RECT  2.8 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.705 ;
      RECT  9.52 -0.14 11.76 0.14 ;
      RECT  9.91 0.14 10.25 0.465 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 1.005 ;
      RECT  1.005 1.005 3.53 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.16 1.565 18.44 1.795 ;
      RECT  15.565 1.795 15.795 3.245 ;
      RECT  15.16 3.245 18.44 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 7.45 0.6 ;
      RECT  11.59 0.37 14.17 0.6 ;
      RECT  7.725 0.695 9.945 0.925 ;
      RECT  7.725 0.925 7.955 1.005 ;
      RECT  9.715 0.925 9.945 1.005 ;
      RECT  6.9 1.005 7.955 1.235 ;
      RECT  9.715 1.005 11.02 1.235 ;
      RECT  12.225 1.005 13.26 1.01 ;
      RECT  12.22 1.01 13.26 1.015 ;
      RECT  12.215 1.015 13.26 1.02 ;
      RECT  12.21 1.02 13.26 1.025 ;
      RECT  12.205 1.025 13.26 1.03 ;
      RECT  12.2 1.03 13.26 1.035 ;
      RECT  12.195 1.035 13.26 1.04 ;
      RECT  12.19 1.04 13.26 1.045 ;
      RECT  12.185 1.045 13.26 1.05 ;
      RECT  12.18 1.05 13.26 1.055 ;
      RECT  12.175 1.055 13.26 1.06 ;
      RECT  12.17 1.06 13.26 1.065 ;
      RECT  12.165 1.065 13.26 1.07 ;
      RECT  12.16 1.07 13.26 1.075 ;
      RECT  12.155 1.075 13.26 1.08 ;
      RECT  12.15 1.08 13.26 1.085 ;
      RECT  12.145 1.085 13.26 1.09 ;
      RECT  12.14 1.09 13.26 1.095 ;
      RECT  12.135 1.095 13.26 1.1 ;
      RECT  12.13 1.1 13.26 1.105 ;
      RECT  12.125 1.105 13.26 1.11 ;
      RECT  12.12 1.11 13.26 1.115 ;
      RECT  12.115 1.115 13.26 1.12 ;
      RECT  12.11 1.12 13.26 1.125 ;
      RECT  12.105 1.125 13.26 1.13 ;
      RECT  12.1 1.13 13.26 1.135 ;
      RECT  12.095 1.135 13.26 1.14 ;
      RECT  12.09 1.14 13.26 1.145 ;
      RECT  12.085 1.145 13.26 1.15 ;
      RECT  12.08 1.15 13.26 1.155 ;
      RECT  12.075 1.155 13.26 1.16 ;
      RECT  12.07 1.16 13.26 1.165 ;
      RECT  12.065 1.165 13.26 1.17 ;
      RECT  12.06 1.17 13.26 1.175 ;
      RECT  12.055 1.175 13.26 1.18 ;
      RECT  12.05 1.18 13.26 1.185 ;
      RECT  12.045 1.185 13.26 1.19 ;
      RECT  12.04 1.19 13.26 1.195 ;
      RECT  12.035 1.195 13.26 1.2 ;
      RECT  12.03 1.2 13.26 1.205 ;
      RECT  12.025 1.205 13.26 1.21 ;
      RECT  12.02 1.21 13.26 1.215 ;
      RECT  12.015 1.215 13.26 1.22 ;
      RECT  12.01 1.22 13.26 1.225 ;
      RECT  12.005 1.225 13.26 1.23 ;
      RECT  12.0 1.23 13.26 1.235 ;
      RECT  11.995 1.235 12.32 1.24 ;
      RECT  11.99 1.24 12.315 1.245 ;
      RECT  11.985 1.245 12.31 1.25 ;
      RECT  11.98 1.25 12.305 1.255 ;
      RECT  11.975 1.255 12.3 1.26 ;
      RECT  11.97 1.26 12.295 1.265 ;
      RECT  11.965 1.265 12.29 1.27 ;
      RECT  11.96 1.27 12.285 1.275 ;
      RECT  11.955 1.275 12.28 1.28 ;
      RECT  11.95 1.28 12.275 1.285 ;
      RECT  11.945 1.285 12.27 1.29 ;
      RECT  11.94 1.29 12.265 1.295 ;
      RECT  11.935 1.295 12.26 1.3 ;
      RECT  11.93 1.3 12.255 1.305 ;
      RECT  11.925 1.305 12.25 1.31 ;
      RECT  11.92 1.31 12.245 1.315 ;
      RECT  11.915 1.315 12.24 1.32 ;
      RECT  11.91 1.32 12.235 1.325 ;
      RECT  11.905 1.325 12.23 1.33 ;
      RECT  11.9 1.33 12.225 1.335 ;
      RECT  11.895 1.335 12.22 1.34 ;
      RECT  11.89 1.34 12.215 1.345 ;
      RECT  11.885 1.345 12.21 1.35 ;
      RECT  11.88 1.35 12.205 1.355 ;
      RECT  11.875 1.355 12.2 1.36 ;
      RECT  11.87 1.36 12.195 1.365 ;
      RECT  11.865 1.365 12.19 1.37 ;
      RECT  11.86 1.37 12.185 1.375 ;
      RECT  11.855 1.375 12.18 1.38 ;
      RECT  11.85 1.38 12.175 1.385 ;
      RECT  11.845 1.385 12.17 1.39 ;
      RECT  11.84 1.39 12.165 1.395 ;
      RECT  11.835 1.395 12.16 1.4 ;
      RECT  11.83 1.4 12.155 1.405 ;
      RECT  11.825 1.405 12.15 1.41 ;
      RECT  11.82 1.41 12.145 1.415 ;
      RECT  11.815 1.415 12.14 1.42 ;
      RECT  11.81 1.42 12.135 1.425 ;
      RECT  11.805 1.425 12.13 1.43 ;
      RECT  11.8 1.43 12.125 1.435 ;
      RECT  11.795 1.435 12.12 1.44 ;
      RECT  11.79 1.44 12.115 1.445 ;
      RECT  11.785 1.445 12.11 1.45 ;
      RECT  11.78 1.45 12.105 1.455 ;
      RECT  11.775 1.455 12.1 1.46 ;
      RECT  11.77 1.46 12.095 1.465 ;
      RECT  11.765 1.465 12.09 1.47 ;
      RECT  11.76 1.47 12.085 1.475 ;
      RECT  11.755 1.475 12.08 1.48 ;
      RECT  11.75 1.48 12.075 1.485 ;
      RECT  11.745 1.485 12.07 1.49 ;
      RECT  11.74 1.49 12.065 1.495 ;
      RECT  11.735 1.495 12.06 1.5 ;
      RECT  11.735 1.5 12.055 1.505 ;
      RECT  11.735 1.505 12.05 1.51 ;
      RECT  11.735 1.51 12.045 1.515 ;
      RECT  11.735 1.515 12.04 1.52 ;
      RECT  11.735 1.52 12.035 1.525 ;
      RECT  11.735 1.525 12.03 1.53 ;
      RECT  11.735 1.53 12.025 1.535 ;
      RECT  11.735 1.535 12.02 1.54 ;
      RECT  11.735 1.54 12.015 1.545 ;
      RECT  11.735 1.545 12.01 1.55 ;
      RECT  11.735 1.55 12.005 1.555 ;
      RECT  11.735 1.555 12.0 1.56 ;
      RECT  11.735 1.56 11.995 1.565 ;
      RECT  11.735 1.565 11.99 1.57 ;
      RECT  11.735 1.57 11.985 1.575 ;
      RECT  11.735 1.575 11.98 1.58 ;
      RECT  11.735 1.58 11.975 1.585 ;
      RECT  11.735 1.585 11.97 1.59 ;
      RECT  11.735 1.59 11.965 3.245 ;
      RECT  11.38 3.245 11.965 3.475 ;
      RECT  11.275 0.89 11.72 1.12 ;
      RECT  11.275 1.12 11.505 1.615 ;
      RECT  7.67 1.615 11.505 1.845 ;
      RECT  8.845 1.845 9.075 3.245 ;
      RECT  7.67 3.245 10.195 3.475 ;
      RECT  9.965 3.475 10.195 3.755 ;
      RECT  9.965 3.755 12.435 3.985 ;
      RECT  12.205 3.985 12.435 4.365 ;
      RECT  12.205 4.365 13.26 4.595 ;
      RECT  3.96 1.005 6.54 1.235 ;
      RECT  8.44 1.155 9.48 1.385 ;
      RECT  0.18 1.565 1.235 1.795 ;
      RECT  1.005 1.795 1.235 4.365 ;
      RECT  0.18 4.365 1.74 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 2.245 4.035 ;
      RECT  2.015 4.035 2.245 4.605 ;
      RECT  2.015 4.605 4.035 4.835 ;
      RECT  3.805 4.835 4.035 5.0 ;
      RECT  3.805 5.0 6.33 5.23 ;
      RECT  2.42 1.565 5.0 1.795 ;
      RECT  13.325 1.565 13.96 1.795 ;
      RECT  13.325 1.795 13.555 2.405 ;
      RECT  12.71 2.405 13.555 2.635 ;
      RECT  13.325 2.635 13.555 3.245 ;
      RECT  13.325 3.245 13.96 3.475 ;
      RECT  5.99 2.405 8.57 2.635 ;
      RECT  5.485 1.51 5.715 3.455 ;
      RECT  2.475 3.685 6.54 3.915 ;
      RECT  6.2 3.915 6.54 4.035 ;
      RECT  2.475 3.915 2.705 4.09 ;
      RECT  6.9 3.705 9.48 3.935 ;
      RECT  6.9 3.935 7.24 3.99 ;
      RECT  3.96 4.145 5.0 4.375 ;
      RECT  8.44 4.215 11.02 4.445 ;
      RECT  16.19 4.405 17.42 4.635 ;
      RECT  16.19 4.635 16.42 5.0 ;
      RECT  17.19 4.635 17.42 5.0 ;
      RECT  12.205 1.695 12.435 3.245 ;
      RECT  12.205 3.245 12.995 3.475 ;
      RECT  12.765 3.475 12.995 3.805 ;
      RECT  12.765 3.805 14.115 4.035 ;
      RECT  13.885 4.035 14.115 4.365 ;
      RECT  13.885 4.365 15.18 4.595 ;
      RECT  14.95 4.595 15.18 5.0 ;
      RECT  14.95 5.0 16.42 5.22 ;
      RECT  17.19 5.0 18.65 5.23 ;
      RECT  14.95 5.22 16.41 5.23 ;
      RECT  5.43 4.48 7.955 4.675 ;
      RECT  5.43 4.675 11.72 4.71 ;
      RECT  11.38 4.48 11.72 4.675 ;
      RECT  7.725 4.71 11.72 4.905 ;
  END
END MDN_MUX4_4
#-----------------------------------------------------------------------
#      Cell        : MDN_MUXI2_3
#      Description : 2-1 multiplexer with inverted output
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUXI2_3
  CLASS CORE ;
  FOREIGN MDN_MUXI2_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.705 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 10.195 1.795 ;
      RECT  9.965 1.795 10.195 3.245 ;
      RECT  6.9 3.245 10.195 3.475 ;
    END
    ANTENNADIFFAREA 4.536 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 4.09 0.6 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.245 1.005 6.22 1.235 ;
      RECT  3.245 1.235 3.475 3.53 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.805 ;
      RECT  1.72 3.805 2.915 4.035 ;
      RECT  3.96 1.565 5.005 1.795 ;
      RECT  6.255 1.51 6.485 2.405 ;
      RECT  6.255 2.405 9.69 2.635 ;
      RECT  6.255 2.635 6.485 3.53 ;
      RECT  3.245 3.805 5.0 4.035 ;
      RECT  3.245 4.035 3.475 4.365 ;
      RECT  2.42 4.365 3.475 4.595 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 4.925 ;
      RECT  0.18 4.365 1.795 4.595 ;
      RECT  1.565 4.595 1.795 4.925 ;
      RECT  1.565 4.925 4.035 5.155 ;
  END
END MDN_MUXI2_3
#-----------------------------------------------------------------------
#      Cell        : MDN_MUXI2_4
#      Description : 2-1 multiplexer with inverted output
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUXI2_4
  CLASS CORE ;
  FOREIGN MDN_MUXI2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.565 11.02 1.795 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  6.9 3.245 11.02 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 4.09 0.6 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.245 1.005 6.22 1.235 ;
      RECT  3.245 1.235 3.475 3.53 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.805 ;
      RECT  1.72 3.805 2.915 4.035 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  6.255 1.51 6.485 2.405 ;
      RECT  6.255 2.405 8.57 2.635 ;
      RECT  6.255 2.635 6.485 3.53 ;
      RECT  9.35 2.405 10.81 2.635 ;
      RECT  3.245 3.805 5.0 4.035 ;
      RECT  3.245 4.035 3.475 4.365 ;
      RECT  2.42 4.365 3.475 4.595 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 4.925 ;
      RECT  0.18 4.365 1.795 4.595 ;
      RECT  1.565 4.595 1.795 4.925 ;
      RECT  1.565 4.925 4.035 5.155 ;
      RECT  8.23 5.0 9.69 5.23 ;
  END
END MDN_MUXI2_4
#-----------------------------------------------------------------------
#      Cell        : MDN_MUXI2_1
#      Description : 2-1 multiplexer with inverted output
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUXI2_1
  CLASS CORE ;
  FOREIGN MDN_MUXI2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  4.31 5.46 5.715 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  0.56 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  4.31 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  1.005 -0.14 1.68 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 1.51 3.475 3.53 ;
    END
    ANTENNADIFFAREA 2.566 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.09 0.445 ;
      RECT  1.565 0.445 4.09 0.675 ;
      RECT  1.565 0.675 1.795 1.565 ;
      RECT  1.565 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 3.245 ;
      RECT  1.72 3.245 2.355 3.475 ;
      RECT  2.42 1.005 5.0 1.235 ;
      RECT  5.485 1.005 6.54 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  3.96 1.565 5.715 1.795 ;
      RECT  4.365 3.805 5.0 4.035 ;
      RECT  4.365 4.035 4.595 4.365 ;
      RECT  3.96 4.365 4.595 4.595 ;
      RECT  4.925 4.365 6.54 4.595 ;
      RECT  4.925 4.595 5.155 4.925 ;
      RECT  2.42 4.365 3.475 4.595 ;
      RECT  3.245 4.595 3.475 4.925 ;
      RECT  3.245 4.925 5.155 5.155 ;
      RECT  1.51 5.0 2.97 5.23 ;
  END
END MDN_MUXI2_1
#-----------------------------------------------------------------------
#      Cell        : MDN_MUXI2_2
#      Description : 2-1 multiplexer with inverted output
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUXI2_2
  CLASS CORE ;
  FOREIGN MDN_MUXI2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 1.82 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 7.42 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.895 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 5.77 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  2.42 3.245 5.77 3.475 ;
    END
    ANTENNADIFFAREA 5.59 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.76 0.37 4.1 0.445 ;
      RECT  3.76 0.445 7.185 0.675 ;
      RECT  6.955 0.675 7.185 1.29 ;
      RECT  8.23 0.37 9.69 0.6 ;
      RECT  2.125 0.445 3.53 0.675 ;
      RECT  2.125 0.675 2.355 1.005 ;
      RECT  0.18 1.005 2.355 1.235 ;
      RECT  7.725 1.005 9.48 1.235 ;
      RECT  7.725 1.235 7.955 1.565 ;
      RECT  4.66 1.005 6.54 1.235 ;
      RECT  6.31 1.235 6.54 1.565 ;
      RECT  6.31 1.565 7.955 1.795 ;
      RECT  2.63 2.405 3.95 2.635 ;
      RECT  3.19 3.805 7.955 4.035 ;
      RECT  7.725 4.035 7.955 4.365 ;
      RECT  7.725 4.365 9.48 4.595 ;
      RECT  3.245 4.365 6.54 4.595 ;
      RECT  3.245 4.595 3.475 4.925 ;
      RECT  0.95 4.925 3.475 5.155 ;
      RECT  6.955 4.31 7.185 4.925 ;
      RECT  3.75 4.925 7.185 5.155 ;
      RECT  3.75 5.155 4.09 5.23 ;
  END
END MDN_MUXI2_2
#-----------------------------------------------------------------------
#      Cell        : MDN_MUXI4_1
#      Description : 4-1 multiplexer with inverted output
#      Equation    : X=!((D0&!S0&!S1)|(D1&S0&!S1)|(D2&!S0&S1)|(D3&S0&S1))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUXI4_1
  CLASS CORE ;
  FOREIGN MDN_MUXI4_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D2
  PIN D3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D3
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 14.14 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.87 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 10.64 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  9.52 -0.14 10.64 0.14 ;
      RECT  9.91 0.14 10.25 0.465 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 1.005 ;
      RECT  1.005 1.005 3.53 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.86 1.565 16.915 1.795 ;
      RECT  16.685 1.795 16.915 3.245 ;
      RECT  15.86 3.245 16.915 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.445 ;
      RECT  1.51 0.445 7.45 0.675 ;
      RECT  4.87 0.37 5.21 0.445 ;
      RECT  7.11 0.37 7.45 0.445 ;
      RECT  11.59 0.37 14.17 0.6 ;
      RECT  7.725 0.745 9.94 0.975 ;
      RECT  7.725 0.975 7.955 1.005 ;
      RECT  9.71 0.975 9.94 1.005 ;
      RECT  6.9 1.005 7.955 1.235 ;
      RECT  9.71 1.005 11.02 1.235 ;
      RECT  12.22 1.005 13.26 1.01 ;
      RECT  12.215 1.01 13.26 1.015 ;
      RECT  12.21 1.015 13.26 1.02 ;
      RECT  12.205 1.02 13.26 1.025 ;
      RECT  12.2 1.025 13.26 1.03 ;
      RECT  12.195 1.03 13.26 1.035 ;
      RECT  12.19 1.035 13.26 1.04 ;
      RECT  12.185 1.04 13.26 1.045 ;
      RECT  12.18 1.045 13.26 1.05 ;
      RECT  12.175 1.05 13.26 1.055 ;
      RECT  12.17 1.055 13.26 1.06 ;
      RECT  12.165 1.06 13.26 1.065 ;
      RECT  12.16 1.065 13.26 1.07 ;
      RECT  12.155 1.07 13.26 1.075 ;
      RECT  12.15 1.075 13.26 1.08 ;
      RECT  12.145 1.08 13.26 1.085 ;
      RECT  12.14 1.085 13.26 1.09 ;
      RECT  12.135 1.09 13.26 1.095 ;
      RECT  12.13 1.095 13.26 1.1 ;
      RECT  12.125 1.1 13.26 1.105 ;
      RECT  12.12 1.105 13.26 1.11 ;
      RECT  12.115 1.11 13.26 1.115 ;
      RECT  12.11 1.115 13.26 1.12 ;
      RECT  12.105 1.12 13.26 1.125 ;
      RECT  12.1 1.125 13.26 1.13 ;
      RECT  12.095 1.13 13.26 1.135 ;
      RECT  12.09 1.135 13.26 1.14 ;
      RECT  12.085 1.14 13.26 1.145 ;
      RECT  12.08 1.145 13.26 1.15 ;
      RECT  12.075 1.15 13.26 1.155 ;
      RECT  12.07 1.155 13.26 1.16 ;
      RECT  12.065 1.16 13.26 1.165 ;
      RECT  12.06 1.165 13.26 1.17 ;
      RECT  12.055 1.17 13.26 1.175 ;
      RECT  12.05 1.175 13.26 1.18 ;
      RECT  12.045 1.18 13.26 1.185 ;
      RECT  12.04 1.185 13.26 1.19 ;
      RECT  12.035 1.19 13.26 1.195 ;
      RECT  12.03 1.195 13.26 1.2 ;
      RECT  12.025 1.2 13.26 1.205 ;
      RECT  12.02 1.205 13.26 1.21 ;
      RECT  12.015 1.21 13.26 1.215 ;
      RECT  12.01 1.215 13.26 1.22 ;
      RECT  12.005 1.22 13.26 1.225 ;
      RECT  12.0 1.225 13.26 1.23 ;
      RECT  11.995 1.23 13.26 1.235 ;
      RECT  11.99 1.235 12.315 1.24 ;
      RECT  11.985 1.24 12.31 1.245 ;
      RECT  11.98 1.245 12.305 1.25 ;
      RECT  11.975 1.25 12.3 1.255 ;
      RECT  11.97 1.255 12.295 1.26 ;
      RECT  11.965 1.26 12.29 1.265 ;
      RECT  11.96 1.265 12.285 1.27 ;
      RECT  11.955 1.27 12.28 1.275 ;
      RECT  11.95 1.275 12.275 1.28 ;
      RECT  11.945 1.28 12.27 1.285 ;
      RECT  11.94 1.285 12.265 1.29 ;
      RECT  11.935 1.29 12.26 1.295 ;
      RECT  11.93 1.295 12.255 1.3 ;
      RECT  11.925 1.3 12.25 1.305 ;
      RECT  11.92 1.305 12.245 1.31 ;
      RECT  11.915 1.31 12.24 1.315 ;
      RECT  11.91 1.315 12.235 1.32 ;
      RECT  11.905 1.32 12.23 1.325 ;
      RECT  11.9 1.325 12.225 1.33 ;
      RECT  11.895 1.33 12.22 1.335 ;
      RECT  11.89 1.335 12.215 1.34 ;
      RECT  11.885 1.34 12.21 1.345 ;
      RECT  11.88 1.345 12.205 1.35 ;
      RECT  11.875 1.35 12.2 1.355 ;
      RECT  11.87 1.355 12.195 1.36 ;
      RECT  11.865 1.36 12.19 1.365 ;
      RECT  11.86 1.365 12.185 1.37 ;
      RECT  11.855 1.37 12.18 1.375 ;
      RECT  11.85 1.375 12.175 1.38 ;
      RECT  11.845 1.38 12.17 1.385 ;
      RECT  11.84 1.385 12.165 1.39 ;
      RECT  11.835 1.39 12.16 1.395 ;
      RECT  11.83 1.395 12.155 1.4 ;
      RECT  11.825 1.4 12.15 1.405 ;
      RECT  11.82 1.405 12.145 1.41 ;
      RECT  11.815 1.41 12.14 1.415 ;
      RECT  11.81 1.415 12.135 1.42 ;
      RECT  11.805 1.42 12.13 1.425 ;
      RECT  11.8 1.425 12.125 1.43 ;
      RECT  11.795 1.43 12.12 1.435 ;
      RECT  11.79 1.435 12.115 1.44 ;
      RECT  11.785 1.44 12.11 1.445 ;
      RECT  11.78 1.445 12.105 1.45 ;
      RECT  11.775 1.45 12.1 1.455 ;
      RECT  11.77 1.455 12.095 1.46 ;
      RECT  11.765 1.46 12.09 1.465 ;
      RECT  11.76 1.465 12.085 1.47 ;
      RECT  11.755 1.47 12.08 1.475 ;
      RECT  11.75 1.475 12.075 1.48 ;
      RECT  11.745 1.48 12.07 1.485 ;
      RECT  11.74 1.485 12.065 1.49 ;
      RECT  11.735 1.49 12.06 1.495 ;
      RECT  11.735 1.495 12.055 1.5 ;
      RECT  11.735 1.5 12.05 1.505 ;
      RECT  11.735 1.505 12.045 1.51 ;
      RECT  11.735 1.51 12.04 1.515 ;
      RECT  11.735 1.515 12.035 1.52 ;
      RECT  11.735 1.52 12.03 1.525 ;
      RECT  11.735 1.525 12.025 1.53 ;
      RECT  11.735 1.53 12.02 1.535 ;
      RECT  11.735 1.535 12.015 1.54 ;
      RECT  11.735 1.54 12.01 1.545 ;
      RECT  11.735 1.545 12.005 1.55 ;
      RECT  11.735 1.55 12.0 1.555 ;
      RECT  11.735 1.555 11.995 1.56 ;
      RECT  11.735 1.56 11.99 1.565 ;
      RECT  11.735 1.565 11.985 1.57 ;
      RECT  11.735 1.57 11.98 1.575 ;
      RECT  11.735 1.575 11.975 1.58 ;
      RECT  11.735 1.58 11.97 1.585 ;
      RECT  11.735 1.585 11.965 3.245 ;
      RECT  11.38 3.245 11.965 3.475 ;
      RECT  11.27 0.89 11.72 1.12 ;
      RECT  11.27 1.12 11.5 1.565 ;
      RECT  9.965 1.565 11.5 1.665 ;
      RECT  7.67 1.665 11.5 1.795 ;
      RECT  7.67 1.795 10.195 1.895 ;
      RECT  8.845 1.895 9.075 3.245 ;
      RECT  7.67 3.245 10.195 3.475 ;
      RECT  9.965 3.475 10.195 3.755 ;
      RECT  9.965 3.755 12.435 3.985 ;
      RECT  12.205 3.985 12.435 4.365 ;
      RECT  12.205 4.365 13.26 4.595 ;
      RECT  3.96 1.005 6.54 1.235 ;
      RECT  8.44 1.205 9.48 1.435 ;
      RECT  0.18 1.565 1.235 1.795 ;
      RECT  1.005 1.795 1.235 4.365 ;
      RECT  0.18 4.365 1.74 4.595 ;
      RECT  1.51 4.595 1.74 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 2.355 4.035 ;
      RECT  2.125 4.035 2.355 4.365 ;
      RECT  2.125 4.365 4.035 4.595 ;
      RECT  3.805 4.595 4.035 5.0 ;
      RECT  3.805 5.0 6.33 5.23 ;
      RECT  2.42 1.565 5.0 1.795 ;
      RECT  13.325 1.565 13.96 1.795 ;
      RECT  13.325 1.795 13.555 2.405 ;
      RECT  12.71 2.405 13.555 2.635 ;
      RECT  13.325 2.635 13.555 3.245 ;
      RECT  13.325 3.245 13.965 3.475 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 2.385 ;
      RECT  15.005 2.385 16.215 2.615 ;
      RECT  15.005 2.615 15.235 3.245 ;
      RECT  15.005 3.245 15.5 3.475 ;
      RECT  5.99 2.415 8.57 2.645 ;
      RECT  12.205 1.695 12.435 3.245 ;
      RECT  12.205 3.245 12.995 3.475 ;
      RECT  12.205 3.475 12.435 3.48 ;
      RECT  12.765 3.475 12.995 3.805 ;
      RECT  12.765 3.805 14.115 4.035 ;
      RECT  13.885 4.035 14.115 4.365 ;
      RECT  13.885 4.365 15.18 4.595 ;
      RECT  14.95 4.595 15.18 5.0 ;
      RECT  14.95 5.0 15.29 5.23 ;
      RECT  2.42 3.245 2.915 3.475 ;
      RECT  2.685 3.475 2.915 3.805 ;
      RECT  2.685 3.805 6.54 4.035 ;
      RECT  3.96 3.245 5.0 3.475 ;
      RECT  5.485 1.59 5.715 3.53 ;
      RECT  6.9 3.755 9.48 3.985 ;
      RECT  8.44 4.215 11.02 4.445 ;
      RECT  5.43 4.54 8.205 4.675 ;
      RECT  5.43 4.675 11.665 4.77 ;
      RECT  11.435 4.425 11.665 4.675 ;
      RECT  7.975 4.77 11.665 4.905 ;
  END
END MDN_MUXI4_1
#-----------------------------------------------------------------------
#      Cell        : MDN_MUXI4_2
#      Description : 4-1 multiplexer with inverted output
#      Equation    : X=!((D0&!S0&!S1)|(D1&S0&!S1)|(D2&!S0&S1)|(D3&S0&S1))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUXI4_2
  CLASS CORE ;
  FOREIGN MDN_MUXI4_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D2
  PIN D3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D3
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 14.14 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.87 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  8.4 5.46 10.64 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  8.4 -0.14 10.64 0.14 ;
      RECT  9.91 0.14 10.25 0.465 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 1.005 ;
      RECT  1.005 1.005 3.53 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.86 1.565 17.74 1.795 ;
      RECT  16.685 1.795 16.915 3.245 ;
      RECT  15.86 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.445 ;
      RECT  1.51 0.445 7.45 0.675 ;
      RECT  4.87 0.37 5.21 0.445 ;
      RECT  7.11 0.37 7.45 0.445 ;
      RECT  11.59 0.37 14.17 0.6 ;
      RECT  17.19 0.37 17.53 0.6 ;
      RECT  17.19 0.6 17.42 1.005 ;
      RECT  16.07 0.37 16.41 0.6 ;
      RECT  16.18 0.6 16.41 1.005 ;
      RECT  16.18 1.005 17.42 1.235 ;
      RECT  7.725 0.695 9.94 0.925 ;
      RECT  7.725 0.925 7.955 1.005 ;
      RECT  9.71 0.925 9.94 1.005 ;
      RECT  6.9 1.005 7.955 1.235 ;
      RECT  9.71 1.005 11.02 1.235 ;
      RECT  12.2 1.005 13.26 1.01 ;
      RECT  12.195 1.01 13.26 1.015 ;
      RECT  12.19 1.015 13.26 1.02 ;
      RECT  12.185 1.02 13.26 1.025 ;
      RECT  12.18 1.025 13.26 1.03 ;
      RECT  12.175 1.03 13.26 1.035 ;
      RECT  12.17 1.035 13.26 1.04 ;
      RECT  12.165 1.04 13.26 1.045 ;
      RECT  12.16 1.045 13.26 1.05 ;
      RECT  12.155 1.05 13.26 1.055 ;
      RECT  12.15 1.055 13.26 1.06 ;
      RECT  12.145 1.06 13.26 1.065 ;
      RECT  12.14 1.065 13.26 1.07 ;
      RECT  12.135 1.07 13.26 1.075 ;
      RECT  12.13 1.075 13.26 1.08 ;
      RECT  12.125 1.08 13.26 1.085 ;
      RECT  12.12 1.085 13.26 1.09 ;
      RECT  12.115 1.09 13.26 1.095 ;
      RECT  12.11 1.095 13.26 1.1 ;
      RECT  12.105 1.1 13.26 1.105 ;
      RECT  12.1 1.105 13.26 1.11 ;
      RECT  12.095 1.11 13.26 1.115 ;
      RECT  12.09 1.115 13.26 1.12 ;
      RECT  12.085 1.12 13.26 1.125 ;
      RECT  12.08 1.125 13.26 1.13 ;
      RECT  12.075 1.13 13.26 1.135 ;
      RECT  12.07 1.135 13.26 1.14 ;
      RECT  12.065 1.14 13.26 1.145 ;
      RECT  12.06 1.145 13.26 1.15 ;
      RECT  12.055 1.15 13.26 1.155 ;
      RECT  12.05 1.155 13.26 1.16 ;
      RECT  12.045 1.16 13.26 1.165 ;
      RECT  12.04 1.165 13.26 1.17 ;
      RECT  12.035 1.17 13.26 1.175 ;
      RECT  12.03 1.175 13.26 1.18 ;
      RECT  12.025 1.18 13.26 1.185 ;
      RECT  12.02 1.185 13.26 1.19 ;
      RECT  12.015 1.19 13.26 1.195 ;
      RECT  12.01 1.195 13.26 1.2 ;
      RECT  12.005 1.2 13.26 1.205 ;
      RECT  12.0 1.205 13.26 1.21 ;
      RECT  11.995 1.21 13.26 1.215 ;
      RECT  11.99 1.215 13.26 1.22 ;
      RECT  11.985 1.22 13.26 1.225 ;
      RECT  11.98 1.225 13.26 1.23 ;
      RECT  11.975 1.23 13.26 1.235 ;
      RECT  11.97 1.235 12.295 1.24 ;
      RECT  11.965 1.24 12.29 1.245 ;
      RECT  11.96 1.245 12.285 1.25 ;
      RECT  11.955 1.25 12.28 1.255 ;
      RECT  11.95 1.255 12.275 1.26 ;
      RECT  11.945 1.26 12.27 1.265 ;
      RECT  11.94 1.265 12.265 1.27 ;
      RECT  11.935 1.27 12.26 1.275 ;
      RECT  11.93 1.275 12.255 1.28 ;
      RECT  11.925 1.28 12.25 1.285 ;
      RECT  11.92 1.285 12.245 1.29 ;
      RECT  11.915 1.29 12.24 1.295 ;
      RECT  11.91 1.295 12.235 1.3 ;
      RECT  11.905 1.3 12.23 1.305 ;
      RECT  11.9 1.305 12.225 1.31 ;
      RECT  11.895 1.31 12.22 1.315 ;
      RECT  11.89 1.315 12.215 1.32 ;
      RECT  11.885 1.32 12.21 1.325 ;
      RECT  11.88 1.325 12.205 1.33 ;
      RECT  11.875 1.33 12.2 1.335 ;
      RECT  11.87 1.335 12.195 1.34 ;
      RECT  11.865 1.34 12.19 1.345 ;
      RECT  11.86 1.345 12.185 1.35 ;
      RECT  11.855 1.35 12.18 1.355 ;
      RECT  11.85 1.355 12.175 1.36 ;
      RECT  11.845 1.36 12.17 1.365 ;
      RECT  11.84 1.365 12.165 1.37 ;
      RECT  11.835 1.37 12.16 1.375 ;
      RECT  11.83 1.375 12.155 1.38 ;
      RECT  11.825 1.38 12.15 1.385 ;
      RECT  11.82 1.385 12.145 1.39 ;
      RECT  11.815 1.39 12.14 1.395 ;
      RECT  11.81 1.395 12.135 1.4 ;
      RECT  11.805 1.4 12.13 1.405 ;
      RECT  11.8 1.405 12.125 1.41 ;
      RECT  11.795 1.41 12.12 1.415 ;
      RECT  11.79 1.415 12.115 1.42 ;
      RECT  11.785 1.42 12.11 1.425 ;
      RECT  11.78 1.425 12.105 1.43 ;
      RECT  11.775 1.43 12.1 1.435 ;
      RECT  11.77 1.435 12.095 1.44 ;
      RECT  11.765 1.44 12.09 1.445 ;
      RECT  11.76 1.445 12.085 1.45 ;
      RECT  11.755 1.45 12.08 1.455 ;
      RECT  11.75 1.455 12.075 1.46 ;
      RECT  11.745 1.46 12.07 1.465 ;
      RECT  11.745 1.465 12.065 1.47 ;
      RECT  11.745 1.47 12.06 1.475 ;
      RECT  11.745 1.475 12.055 1.48 ;
      RECT  11.745 1.48 12.05 1.485 ;
      RECT  11.745 1.485 12.045 1.49 ;
      RECT  11.745 1.49 12.04 1.495 ;
      RECT  11.745 1.495 12.035 1.5 ;
      RECT  11.745 1.5 12.03 1.505 ;
      RECT  11.745 1.505 12.025 1.51 ;
      RECT  11.745 1.51 12.02 1.515 ;
      RECT  11.745 1.515 12.015 1.52 ;
      RECT  11.745 1.52 12.01 1.525 ;
      RECT  11.745 1.525 12.005 1.53 ;
      RECT  11.745 1.53 12.0 1.535 ;
      RECT  11.745 1.535 11.995 1.54 ;
      RECT  11.745 1.54 11.99 1.545 ;
      RECT  11.745 1.545 11.985 1.55 ;
      RECT  11.745 1.55 11.98 1.555 ;
      RECT  11.745 1.555 11.975 3.245 ;
      RECT  11.38 3.245 11.975 3.475 ;
      RECT  11.25 0.89 11.72 1.12 ;
      RECT  11.25 1.12 11.48 1.565 ;
      RECT  9.965 1.565 11.48 1.665 ;
      RECT  7.67 1.665 11.48 1.795 ;
      RECT  7.67 1.795 10.195 1.895 ;
      RECT  8.845 1.895 9.075 3.245 ;
      RECT  7.67 3.245 10.195 3.475 ;
      RECT  9.965 3.475 10.195 3.755 ;
      RECT  9.965 3.755 12.435 3.985 ;
      RECT  12.205 3.985 12.435 4.365 ;
      RECT  12.205 4.365 13.26 4.595 ;
      RECT  3.96 1.005 6.54 1.235 ;
      RECT  8.44 1.17 9.48 1.4 ;
      RECT  0.18 1.565 1.235 1.795 ;
      RECT  1.005 1.795 1.235 4.365 ;
      RECT  0.18 4.365 1.695 4.595 ;
      RECT  1.465 4.595 1.695 5.0 ;
      RECT  1.465 5.0 1.85 5.23 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 2.155 4.035 ;
      RECT  1.925 4.035 2.155 4.365 ;
      RECT  1.925 4.365 4.595 4.595 ;
      RECT  4.365 4.595 4.595 5.0 ;
      RECT  4.365 5.0 6.33 5.23 ;
      RECT  2.42 1.565 5.0 1.795 ;
      RECT  13.325 1.565 13.96 1.795 ;
      RECT  13.325 1.795 13.555 2.405 ;
      RECT  12.71 2.405 13.555 2.635 ;
      RECT  13.325 2.635 13.555 3.245 ;
      RECT  13.325 3.245 13.96 3.475 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 2.395 ;
      RECT  15.005 2.395 16.41 2.625 ;
      RECT  15.005 2.625 15.235 3.245 ;
      RECT  15.005 3.245 15.5 3.475 ;
      RECT  5.99 2.405 8.57 2.635 ;
      RECT  12.205 1.695 12.435 3.245 ;
      RECT  12.205 3.245 12.995 3.475 ;
      RECT  12.765 3.475 12.995 3.805 ;
      RECT  12.765 3.805 15.18 4.035 ;
      RECT  14.95 4.035 15.18 5.0 ;
      RECT  14.95 5.0 15.29 5.23 ;
      RECT  3.96 3.245 5.0 3.475 ;
      RECT  5.485 1.51 5.715 3.53 ;
      RECT  6.9 3.755 9.48 3.985 ;
      RECT  2.42 3.805 6.54 4.035 ;
      RECT  8.44 4.215 11.02 4.445 ;
      RECT  5.43 4.48 7.955 4.675 ;
      RECT  5.43 4.675 11.665 4.71 ;
      RECT  11.435 4.425 11.665 4.675 ;
      RECT  7.725 4.71 11.665 4.905 ;
  END
END MDN_MUXI4_2
#-----------------------------------------------------------------------
#      Cell        : MDN_MUXI4_4
#      Description : 4-1 multiplexer with inverted output
#      Equation    : X=!((D0&!S0&!S1)|(D1&S0&!S1)|(D2&!S0&S1)|(D3&S0&S1))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_MUXI4_4
  CLASS CORE ;
  FOREIGN MDN_MUXI4_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D2
  PIN D3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D3
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 14.14 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  8.4 5.46 10.64 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  8.4 -0.14 10.64 0.14 ;
      RECT  9.91 0.14 10.25 0.465 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 1.005 ;
      RECT  1.005 1.005 3.53 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  15.86 1.565 19.98 1.795 ;
      RECT  17.805 1.795 18.035 3.245 ;
      RECT  15.86 3.245 19.98 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.51 0.37 1.85 0.445 ;
      RECT  1.51 0.445 7.45 0.675 ;
      RECT  4.87 0.37 5.21 0.445 ;
      RECT  7.11 0.37 7.45 0.445 ;
      RECT  11.59 0.37 14.17 0.6 ;
      RECT  17.19 0.37 18.65 0.6 ;
      RECT  7.725 0.695 10.195 0.925 ;
      RECT  7.725 0.925 7.955 1.005 ;
      RECT  9.965 0.925 10.195 1.005 ;
      RECT  6.9 1.005 7.955 1.235 ;
      RECT  9.965 1.005 11.02 1.235 ;
      RECT  12.195 1.005 13.26 1.01 ;
      RECT  12.19 1.01 13.26 1.015 ;
      RECT  12.185 1.015 13.26 1.02 ;
      RECT  12.18 1.02 13.26 1.025 ;
      RECT  12.175 1.025 13.26 1.03 ;
      RECT  12.17 1.03 13.26 1.035 ;
      RECT  12.165 1.035 13.26 1.04 ;
      RECT  12.16 1.04 13.26 1.045 ;
      RECT  12.155 1.045 13.26 1.05 ;
      RECT  12.15 1.05 13.26 1.055 ;
      RECT  12.145 1.055 13.26 1.06 ;
      RECT  12.14 1.06 13.26 1.065 ;
      RECT  12.135 1.065 13.26 1.07 ;
      RECT  12.13 1.07 13.26 1.075 ;
      RECT  12.125 1.075 13.26 1.08 ;
      RECT  12.12 1.08 13.26 1.085 ;
      RECT  12.115 1.085 13.26 1.09 ;
      RECT  12.11 1.09 13.26 1.095 ;
      RECT  12.105 1.095 13.26 1.1 ;
      RECT  12.1 1.1 13.26 1.105 ;
      RECT  12.095 1.105 13.26 1.11 ;
      RECT  12.09 1.11 13.26 1.115 ;
      RECT  12.085 1.115 13.26 1.12 ;
      RECT  12.08 1.12 13.26 1.125 ;
      RECT  12.075 1.125 13.26 1.13 ;
      RECT  12.07 1.13 13.26 1.135 ;
      RECT  12.065 1.135 13.26 1.14 ;
      RECT  12.06 1.14 13.26 1.145 ;
      RECT  12.055 1.145 13.26 1.15 ;
      RECT  12.05 1.15 13.26 1.155 ;
      RECT  12.045 1.155 13.26 1.16 ;
      RECT  12.04 1.16 13.26 1.165 ;
      RECT  12.035 1.165 13.26 1.17 ;
      RECT  12.03 1.17 13.26 1.175 ;
      RECT  12.025 1.175 13.26 1.18 ;
      RECT  12.02 1.18 13.26 1.185 ;
      RECT  12.015 1.185 13.26 1.19 ;
      RECT  12.01 1.19 13.26 1.195 ;
      RECT  12.005 1.195 13.26 1.2 ;
      RECT  12.0 1.2 13.26 1.205 ;
      RECT  11.995 1.205 13.26 1.21 ;
      RECT  11.99 1.21 13.26 1.215 ;
      RECT  11.985 1.215 13.26 1.22 ;
      RECT  11.98 1.22 13.26 1.225 ;
      RECT  11.975 1.225 13.26 1.23 ;
      RECT  11.97 1.23 13.26 1.235 ;
      RECT  11.965 1.235 12.29 1.24 ;
      RECT  11.96 1.24 12.285 1.245 ;
      RECT  11.955 1.245 12.28 1.25 ;
      RECT  11.95 1.25 12.275 1.255 ;
      RECT  11.945 1.255 12.27 1.26 ;
      RECT  11.94 1.26 12.265 1.265 ;
      RECT  11.935 1.265 12.26 1.27 ;
      RECT  11.93 1.27 12.255 1.275 ;
      RECT  11.925 1.275 12.25 1.28 ;
      RECT  11.92 1.28 12.245 1.285 ;
      RECT  11.915 1.285 12.24 1.29 ;
      RECT  11.91 1.29 12.235 1.295 ;
      RECT  11.905 1.295 12.23 1.3 ;
      RECT  11.9 1.3 12.225 1.305 ;
      RECT  11.895 1.305 12.22 1.31 ;
      RECT  11.89 1.31 12.215 1.315 ;
      RECT  11.885 1.315 12.21 1.32 ;
      RECT  11.88 1.32 12.205 1.325 ;
      RECT  11.875 1.325 12.2 1.33 ;
      RECT  11.87 1.33 12.195 1.335 ;
      RECT  11.865 1.335 12.19 1.34 ;
      RECT  11.86 1.34 12.185 1.345 ;
      RECT  11.855 1.345 12.18 1.35 ;
      RECT  11.85 1.35 12.175 1.355 ;
      RECT  11.845 1.355 12.17 1.36 ;
      RECT  11.84 1.36 12.165 1.365 ;
      RECT  11.835 1.365 12.16 1.37 ;
      RECT  11.83 1.37 12.155 1.375 ;
      RECT  11.825 1.375 12.15 1.38 ;
      RECT  11.82 1.38 12.145 1.385 ;
      RECT  11.815 1.385 12.14 1.39 ;
      RECT  11.81 1.39 12.135 1.395 ;
      RECT  11.805 1.395 12.13 1.4 ;
      RECT  11.8 1.4 12.125 1.405 ;
      RECT  11.795 1.405 12.12 1.41 ;
      RECT  11.79 1.41 12.115 1.415 ;
      RECT  11.785 1.415 12.11 1.42 ;
      RECT  11.78 1.42 12.105 1.425 ;
      RECT  11.775 1.425 12.1 1.43 ;
      RECT  11.77 1.43 12.095 1.435 ;
      RECT  11.765 1.435 12.09 1.44 ;
      RECT  11.76 1.44 12.085 1.445 ;
      RECT  11.755 1.445 12.08 1.45 ;
      RECT  11.75 1.45 12.075 1.455 ;
      RECT  11.745 1.455 12.07 1.46 ;
      RECT  11.745 1.46 12.065 1.465 ;
      RECT  11.745 1.465 12.06 1.47 ;
      RECT  11.745 1.47 12.055 1.475 ;
      RECT  11.745 1.475 12.05 1.48 ;
      RECT  11.745 1.48 12.045 1.485 ;
      RECT  11.745 1.485 12.04 1.49 ;
      RECT  11.745 1.49 12.035 1.495 ;
      RECT  11.745 1.495 12.03 1.5 ;
      RECT  11.745 1.5 12.025 1.505 ;
      RECT  11.745 1.505 12.02 1.51 ;
      RECT  11.745 1.51 12.015 1.515 ;
      RECT  11.745 1.515 12.01 1.52 ;
      RECT  11.745 1.52 12.005 1.525 ;
      RECT  11.745 1.525 12.0 1.53 ;
      RECT  11.745 1.53 11.995 1.535 ;
      RECT  11.745 1.535 11.99 1.54 ;
      RECT  11.745 1.54 11.985 1.545 ;
      RECT  11.745 1.545 11.98 1.55 ;
      RECT  11.745 1.55 11.975 3.245 ;
      RECT  11.38 3.245 11.975 3.475 ;
      RECT  11.275 0.89 11.72 1.12 ;
      RECT  11.275 1.12 11.505 1.565 ;
      RECT  9.965 1.565 11.505 1.665 ;
      RECT  7.67 1.665 11.505 1.795 ;
      RECT  7.67 1.795 10.195 1.895 ;
      RECT  8.845 1.895 9.075 3.245 ;
      RECT  7.67 3.245 10.195 3.475 ;
      RECT  9.965 3.475 10.195 3.755 ;
      RECT  9.965 3.755 12.435 3.985 ;
      RECT  12.205 3.985 12.435 4.365 ;
      RECT  12.205 4.365 13.26 4.595 ;
      RECT  3.96 1.005 6.54 1.235 ;
      RECT  8.44 1.155 9.48 1.385 ;
      RECT  0.18 1.565 1.235 1.795 ;
      RECT  1.005 1.795 1.235 4.365 ;
      RECT  0.18 4.365 1.725 4.595 ;
      RECT  1.495 4.595 1.725 5.0 ;
      RECT  1.495 5.0 1.85 5.23 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 3.805 ;
      RECT  1.565 3.805 2.19 4.035 ;
      RECT  1.96 4.035 2.19 4.365 ;
      RECT  1.96 4.365 4.035 4.595 ;
      RECT  3.805 4.595 4.035 5.0 ;
      RECT  3.805 5.0 6.33 5.23 ;
      RECT  2.42 1.565 5.0 1.795 ;
      RECT  13.325 1.565 13.96 1.795 ;
      RECT  13.325 1.795 13.555 2.405 ;
      RECT  12.71 2.405 13.555 2.635 ;
      RECT  13.325 2.635 13.555 3.245 ;
      RECT  13.325 3.245 13.96 3.475 ;
      RECT  15.005 1.565 15.5 1.795 ;
      RECT  15.005 1.795 15.235 2.405 ;
      RECT  15.005 2.405 17.53 2.635 ;
      RECT  15.005 2.635 15.235 3.245 ;
      RECT  15.005 3.245 15.5 3.475 ;
      RECT  5.99 2.405 8.57 2.635 ;
      RECT  18.31 2.405 19.77 2.635 ;
      RECT  12.205 1.695 12.435 3.245 ;
      RECT  12.205 3.245 12.995 3.475 ;
      RECT  12.765 3.475 12.995 3.805 ;
      RECT  12.765 3.805 15.18 4.035 ;
      RECT  14.95 4.035 15.18 5.0 ;
      RECT  14.95 5.0 15.29 5.23 ;
      RECT  3.96 3.245 5.0 3.475 ;
      RECT  5.485 1.51 5.715 3.53 ;
      RECT  6.9 3.755 9.48 3.985 ;
      RECT  2.42 3.805 6.54 4.035 ;
      RECT  8.44 4.215 11.02 4.445 ;
      RECT  5.43 4.365 7.955 4.595 ;
      RECT  7.725 4.595 7.955 4.675 ;
      RECT  7.725 4.675 11.665 4.905 ;
      RECT  11.435 4.425 11.665 4.675 ;
  END
END MDN_MUXI4_4
#-----------------------------------------------------------------------
#      Cell        : MDN_ND2_1
#      Description : 2-Input NAND
#      Equation    : X=!(A1&A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND2_1
  CLASS CORE ;
  FOREIGN MDN_ND2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.24 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.565 4.365 2.06 4.595 ;
      RECT  1.565 4.595 1.795 5.46 ;
      RECT  1.565 5.46 2.41 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 2.24 5.74 ;
      LAYER VIA12 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 2.24 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 1.005 2.06 1.235 ;
      RECT  1.005 1.235 1.235 3.53 ;
    END
    ANTENNADIFFAREA 2.086 ;
  END X
END MDN_ND2_1
#-----------------------------------------------------------------------
#      Cell        : MDN_ND2_12
#      Description : 2-Input NAND
#      Equation    : X=!(A1&A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND2_12
  CLASS CORE ;
  FOREIGN MDN_ND2_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 26.88 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 26.46 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
      RECT  18.34 2.355 18.62 2.915 ;
      RECT  19.46 2.355 19.74 2.915 ;
      RECT  20.58 2.355 20.86 2.915 ;
      RECT  21.7 2.355 21.98 2.915 ;
      RECT  22.82 2.355 23.1 2.915 ;
      RECT  23.94 2.355 24.22 2.915 ;
      RECT  25.06 2.355 25.34 2.915 ;
      RECT  26.18 2.355 26.46 2.915 ;
    END
    ANTENNAGATEAREA 6.804 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 13.02 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 6.804 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 4.905 25.875 5.46 ;
      RECT  25.645 5.46 27.05 5.74 ;
      RECT  23.405 4.905 23.635 5.46 ;
      RECT  22.96 5.46 23.635 5.74 ;
      RECT  21.165 4.905 21.395 5.46 ;
      RECT  21.165 5.46 21.84 5.74 ;
      RECT  18.925 4.905 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  16.685 4.905 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  12.205 4.905 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 4.905 14.675 5.46 ;
      RECT  9.965 4.905 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.905 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.905 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.905 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.905 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 26.88 5.74 ;
      LAYER VIA12 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  26.32 -0.14 27.05 0.14 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.695 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.695 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.695 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.695 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.695 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 26.88 0.14 ;
      LAYER VIA12 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.49 0.985 26.645 1.49 ;
      RECT  13.25 1.49 26.645 1.545 ;
      RECT  13.25 1.545 13.87 1.87 ;
      RECT  13.25 1.87 13.63 4.06 ;
      RECT  0.235 4.06 26.645 4.62 ;
    END
    ANTENNADIFFAREA 28.92 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  13.03 0.445 25.93 0.675 ;
      RECT  13.03 0.675 13.26 1.005 ;
      RECT  0.18 1.005 13.26 1.235 ;
  END
END MDN_ND2_12
#-----------------------------------------------------------------------
#      Cell        : MDN_ND2_16
#      Description : 2-Input NAND
#      Equation    : X=!(A1&A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND2_16
  CLASS CORE ;
  FOREIGN MDN_ND2_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 35.84 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.34 4.365 35.42 4.595 ;
      RECT  18.34 4.595 18.62 5.0 ;
      RECT  19.46 4.595 19.74 5.0 ;
      RECT  20.58 4.595 20.86 5.0 ;
      RECT  21.7 4.595 21.98 5.0 ;
      RECT  22.82 4.595 23.1 5.0 ;
      RECT  23.94 4.595 24.22 5.0 ;
      RECT  25.06 4.595 25.34 5.0 ;
      RECT  26.18 4.595 26.46 5.0 ;
      RECT  27.3 4.595 27.58 5.0 ;
      RECT  28.42 4.595 28.7 5.0 ;
      RECT  29.54 4.595 29.82 5.0 ;
      RECT  30.66 4.595 30.94 5.0 ;
      RECT  31.78 4.595 32.06 5.0 ;
      RECT  32.9 4.595 33.18 5.0 ;
      RECT  34.02 4.595 34.3 5.0 ;
      RECT  35.14 4.595 35.42 5.0 ;
      RECT  18.31 5.0 18.65 5.23 ;
      RECT  19.43 5.0 19.77 5.23 ;
      RECT  20.55 5.0 20.89 5.23 ;
      RECT  21.67 5.0 22.01 5.23 ;
      RECT  22.79 5.0 23.13 5.23 ;
      RECT  23.91 5.0 24.25 5.23 ;
      RECT  25.03 5.0 25.37 5.23 ;
      RECT  26.15 5.0 26.49 5.23 ;
      RECT  27.27 5.0 27.61 5.23 ;
      RECT  28.39 5.0 28.73 5.23 ;
      RECT  29.51 5.0 29.85 5.23 ;
      RECT  30.63 5.0 30.97 5.23 ;
      RECT  31.75 5.0 32.09 5.23 ;
      RECT  32.87 5.0 33.21 5.23 ;
      RECT  33.99 5.0 34.33 5.23 ;
      RECT  35.11 5.0 35.45 5.23 ;
    END
    ANTENNAGATEAREA 9.072 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 17.5 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 9.072 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  34.605 5.08 34.835 5.46 ;
      RECT  34.605 5.46 36.01 5.74 ;
      RECT  32.365 5.08 32.595 5.46 ;
      RECT  32.365 5.46 33.04 5.74 ;
      RECT  30.125 5.08 30.355 5.46 ;
      RECT  30.125 5.46 30.8 5.74 ;
      RECT  27.885 5.08 28.115 5.46 ;
      RECT  27.885 5.46 28.56 5.74 ;
      RECT  25.645 5.08 25.875 5.46 ;
      RECT  25.645 5.46 26.32 5.74 ;
      RECT  23.405 5.08 23.635 5.46 ;
      RECT  23.405 5.46 24.08 5.74 ;
      RECT  21.165 5.08 21.395 5.46 ;
      RECT  21.165 5.46 21.84 5.74 ;
      RECT  16.685 5.08 16.915 5.46 ;
      RECT  16.685 5.46 19.155 5.74 ;
      RECT  18.925 5.08 19.155 5.46 ;
      RECT  14.445 5.08 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  12.205 5.08 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  9.965 5.08 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 5.08 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 5.08 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 5.08 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.565 4.48 2.06 4.71 ;
      RECT  1.565 4.71 1.795 5.46 ;
      RECT  1.565 5.46 2.24 5.74 ;
      RECT  0.18 4.48 0.675 4.71 ;
      RECT  0.445 4.71 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 35.84 5.74 ;
      LAYER VIA12 ;
      RECT  34.87 5.47 35.13 5.73 ;
      RECT  35.43 5.47 35.69 5.73 ;
      RECT  32.63 5.47 32.89 5.73 ;
      RECT  30.39 5.47 30.65 5.73 ;
      RECT  28.15 5.47 28.41 5.73 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  18.07 5.47 18.33 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  35.28 -0.14 36.01 0.14 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.52 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.52 ;
      RECT  11.76 -0.14 12.435 0.14 ;
      RECT  12.205 0.14 12.435 0.52 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.52 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.52 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.52 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.52 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.52 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 35.84 0.14 ;
      LAYER VIA12 ;
      RECT  35.43 -0.13 35.69 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.02 1.54 18.85 1.63 ;
      RECT  18.02 1.63 35.605 2.1 ;
      RECT  18.02 2.1 18.85 2.94 ;
      RECT  26.4 2.1 27.23 2.94 ;
      RECT  34.62 2.1 35.09 2.94 ;
      RECT  18.02 2.94 35.605 3.22 ;
      RECT  17.225 3.22 35.605 3.41 ;
      RECT  17.225 3.41 18.62 3.78 ;
      RECT  0.95 3.78 18.62 4.06 ;
      RECT  0.95 4.06 17.92 4.25 ;
      RECT  2.29 4.25 17.92 4.61 ;
    END
    ANTENNADIFFAREA 38.236 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  17.455 0.445 34.89 0.675 ;
      RECT  17.455 0.675 17.685 1.005 ;
      RECT  0.18 1.005 17.685 1.235 ;
  END
END MDN_ND2_16
#-----------------------------------------------------------------------
#      Cell        : MDN_ND2_2
#      Description : 2-Input NAND
#      Equation    : X=!(A1&A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND2_2
  CLASS CORE ;
  FOREIGN MDN_ND2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.685 ;
      RECT  2.66 2.685 4.06 2.915 ;
      RECT  3.78 2.125 4.06 2.685 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 1.82 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 4.65 5.74 ;
      RECT  1.72 4.365 2.76 4.595 ;
      RECT  2.125 4.595 2.355 5.46 ;
      RECT  1.68 5.46 2.8 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 2.06 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.125 1.565 3.53 1.795 ;
      RECT  2.125 1.795 2.355 3.245 ;
      RECT  0.945 3.245 3.53 3.475 ;
    END
    ANTENNADIFFAREA 4.038 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 2.65 0.675 ;
      RECT  2.42 0.675 2.65 1.005 ;
      RECT  2.42 1.005 4.3 1.235 ;
  END
END MDN_ND2_2
#-----------------------------------------------------------------------
#      Cell        : MDN_ND2_3
#      Description : 2-Input NAND
#      Equation    : X=!(A1&A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND2_3
  CLASS CORE ;
  FOREIGN MDN_ND2_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 6.3 2.355 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.93 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 2.76 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 1.005 6.54 1.235 ;
      RECT  3.245 1.235 3.475 3.805 ;
      RECT  0.18 3.805 6.54 4.035 ;
    END
    ANTENNADIFFAREA 7.23 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 5.77 0.675 ;
  END
END MDN_ND2_3
#-----------------------------------------------------------------------
#      Cell        : MDN_ND2_4
#      Description : 2-Input NAND
#      Equation    : X=!(A1&A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND2_4
  CLASS CORE ;
  FOREIGN MDN_ND2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.695 ;
      RECT  4.9 2.695 8.54 2.915 ;
      RECT  6.02 2.125 6.3 2.695 ;
      RECT  7.14 2.125 7.42 2.695 ;
      RECT  8.26 2.125 8.54 2.695 ;
      RECT  4.925 2.915 8.515 2.925 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.695 ;
      RECT  0.42 2.695 4.06 2.915 ;
      RECT  1.54 2.125 1.82 2.695 ;
      RECT  2.66 2.125 2.94 2.695 ;
      RECT  3.78 2.125 4.06 2.695 ;
      RECT  0.465 2.915 4.035 2.925 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  8.285 4.365 8.78 4.595 ;
      RECT  8.285 4.595 8.515 5.46 ;
      RECT  8.285 5.46 9.13 5.74 ;
      RECT  6.2 4.365 7.24 4.595 ;
      RECT  6.605 4.595 6.835 5.46 ;
      RECT  6.16 5.46 7.28 5.74 ;
      RECT  3.96 4.365 5.0 4.595 ;
      RECT  4.365 4.595 4.595 5.46 ;
      RECT  3.92 5.46 5.04 5.74 ;
      RECT  1.72 4.365 2.76 4.595 ;
      RECT  2.125 4.595 2.355 5.46 ;
      RECT  1.68 5.46 2.8 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      RECT  3.245 0.14 3.475 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.32 1.565 8.01 1.795 ;
      RECT  4.32 1.795 4.85 1.82 ;
      RECT  4.32 1.82 4.64 3.22 ;
      RECT  0.91 3.22 4.85 3.245 ;
      RECT  0.91 3.245 8.01 3.475 ;
      RECT  0.91 3.475 4.85 3.5 ;
    END
    ANTENNADIFFAREA 8.076 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 8.78 1.235 ;
  END
END MDN_ND2_4
#-----------------------------------------------------------------------
#      Cell        : MDN_ND2_6
#      Description : 2-Input NAND
#      Equation    : X=!(A1&A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND2_6
  CLASS CORE ;
  FOREIGN MDN_ND2_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 13.02 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 6.3 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.32 -0.14 13.61 0.14 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 0.98 13.26 1.26 ;
      RECT  7.14 1.26 7.42 1.54 ;
      RECT  6.58 1.54 7.42 1.82 ;
      RECT  6.58 1.82 6.86 3.78 ;
      RECT  0.18 3.78 13.26 4.06 ;
    END
    ANTENNADIFFAREA 14.46 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  6.26 0.42 12.515 0.7 ;
      RECT  6.26 0.7 6.54 0.98 ;
      RECT  0.18 0.98 6.54 1.26 ;
  END
END MDN_ND2_6
#-----------------------------------------------------------------------
#      Cell        : MDN_ND2_8
#      Description : 2-Input NAND
#      Equation    : X=!(A1&A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND2_8
  CLASS CORE ;
  FOREIGN MDN_ND2_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 17.5 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 4.536 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 8.54 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 4.536 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  17.36 -0.14 18.09 0.14 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.335 0.935 17.74 1.305 ;
      RECT  9.335 1.305 9.705 1.495 ;
      RECT  8.77 1.495 9.705 1.865 ;
      RECT  8.77 1.865 9.15 3.735 ;
      RECT  0.18 3.735 17.74 4.105 ;
    END
    ANTENNADIFFAREA 19.28 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.5 0.42 16.97 0.7 ;
      RECT  8.5 0.7 8.78 0.98 ;
      RECT  0.18 0.98 8.78 1.26 ;
  END
END MDN_ND2_8
#-----------------------------------------------------------------------
#      Cell        : MDN_ND2B_1
#      Description : 2-Input NAND (A inverted input)
#      Equation    : X=!(!A&B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND2B_1
  CLASS CORE ;
  FOREIGN MDN_ND2B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 -0.14 4.65 0.14 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  1.005 -0.14 1.68 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 3.805 ;
      RECT  2.42 3.805 4.3 4.035 ;
    END
    ANTENNADIFFAREA 2.41 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
  END
END MDN_ND2B_1
#-----------------------------------------------------------------------
#      Cell        : MDN_ND2B_2
#      Description : 2-Input NAND (A inverted input)
#      Equation    : X=!(!A&B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND2B_2
  CLASS CORE ;
  FOREIGN MDN_ND2B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 -0.14 6.89 0.14 ;
      RECT  6.045 0.14 6.275 1.005 ;
      RECT  4.66 1.005 6.54 1.235 ;
      RECT  1.005 -0.14 1.68 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  3.245 1.565 4.595 1.795 ;
      RECT  4.365 1.795 4.595 3.805 ;
      RECT  2.42 3.805 6.54 4.035 ;
    END
    ANTENNADIFFAREA 4.82 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.445 5.77 0.675 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 2.685 ;
      RECT  2.685 2.685 4.035 2.915 ;
      RECT  3.805 2.35 4.035 2.685 ;
      RECT  2.685 2.915 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
  END
END MDN_ND2B_2
#-----------------------------------------------------------------------
#      Cell        : MDN_ND2B_3
#      Description : 2-Input NAND (A inverted input)
#      Equation    : X=!(!A&B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND2B_3
  CLASS CORE ;
  FOREIGN MDN_ND2B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 8.54 2.355 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  1.005 5.46 2.41 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  8.285 -0.14 9.13 0.14 ;
      RECT  8.285 0.14 8.515 1.005 ;
      RECT  6.2 1.005 8.78 1.235 ;
      RECT  1.005 -0.14 1.68 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 5.715 1.235 ;
      RECT  5.485 1.235 5.715 3.805 ;
      RECT  2.42 3.805 8.78 4.035 ;
    END
    ANTENNADIFFAREA 7.23 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.445 8.01 0.675 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 2.685 ;
      RECT  2.685 2.685 5.155 2.915 ;
      RECT  3.805 2.35 4.035 2.685 ;
      RECT  4.925 2.35 5.155 2.685 ;
      RECT  2.685 2.915 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
  END
END MDN_ND2B_3
#-----------------------------------------------------------------------
#      Cell        : MDN_ND2B_4
#      Description : 2-Input NAND (A inverted input)
#      Equation    : X=!(!A&B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND2B_4
  CLASS CORE ;
  FOREIGN MDN_ND2B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 10.78 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 5.715 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  5.485 1.565 6.835 1.795 ;
      RECT  6.605 1.795 6.835 3.805 ;
      RECT  2.42 3.805 11.02 4.035 ;
    END
    ANTENNADIFFAREA 9.64 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.445 6.835 0.675 ;
      RECT  6.605 0.675 6.835 1.005 ;
      RECT  6.605 1.005 11.02 1.235 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 2.685 ;
      RECT  2.685 2.685 6.275 2.915 ;
      RECT  3.805 2.35 4.035 2.685 ;
      RECT  4.925 2.35 5.155 2.685 ;
      RECT  6.045 2.35 6.275 2.685 ;
      RECT  2.685 2.915 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
  END
END MDN_ND2B_4
#-----------------------------------------------------------------------
#      Cell        : MDN_ND2B_6
#      Description : 2-Input NAND (A inverted input)
#      Equation    : X=!(!A&B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND2B_6
  CLASS CORE ;
  FOREIGN MDN_ND2B_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 1.82 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 15.26 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.565 4.365 2.06 4.595 ;
      RECT  1.565 4.595 1.795 5.46 ;
      RECT  1.565 5.46 2.41 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  11.76 -0.14 12.435 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  1.565 -0.14 2.41 0.14 ;
      RECT  1.565 0.14 1.795 1.005 ;
      RECT  1.565 1.005 2.06 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 0.98 8.54 1.26 ;
      RECT  8.26 1.26 8.54 1.54 ;
      RECT  8.26 1.54 9.1 1.82 ;
      RECT  8.82 1.82 9.1 3.78 ;
      RECT  2.42 3.78 15.5 4.06 ;
    END
    ANTENNADIFFAREA 14.46 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.42 9.1 0.7 ;
      RECT  8.82 0.7 9.1 0.98 ;
      RECT  8.82 0.98 15.5 1.26 ;
      RECT  0.95 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 2.685 ;
      RECT  2.125 2.685 8.515 2.915 ;
      RECT  2.685 2.35 2.915 2.685 ;
      RECT  3.805 2.35 4.035 2.685 ;
      RECT  4.925 2.35 5.155 2.685 ;
      RECT  6.045 2.35 6.275 2.685 ;
      RECT  7.165 2.35 7.395 2.685 ;
      RECT  8.285 2.35 8.515 2.685 ;
      RECT  2.125 2.915 2.355 3.245 ;
      RECT  0.945 3.245 2.355 3.475 ;
  END
END MDN_ND2B_6
#-----------------------------------------------------------------------
#      Cell        : MDN_ND3_1
#      Description : 3-Input NAND
#      Equation    : X=!(A1&A2&A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND3_1
  CLASS CORE ;
  FOREIGN MDN_ND3_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 4.65 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  1.005 5.46 1.68 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 -0.14 2.41 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 1.005 4.3 1.235 ;
      RECT  3.245 1.235 3.475 3.805 ;
      RECT  1.72 3.805 4.3 4.035 ;
    END
    ANTENNADIFFAREA 3.308 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.005 2.76 1.235 ;
  END
END MDN_ND3_1
#-----------------------------------------------------------------------
#      Cell        : MDN_ND3_2
#      Description : 3-Input NAND
#      Equation    : X=!(A1&A2&A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND3_2
  CLASS CORE ;
  FOREIGN MDN_ND3_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.925 1.005 6.54 1.235 ;
      RECT  4.925 1.235 5.155 1.565 ;
      RECT  4.365 1.565 5.155 1.795 ;
      RECT  4.365 1.795 4.595 3.805 ;
      RECT  0.18 3.805 6.54 4.035 ;
    END
    ANTENNADIFFAREA 6.616 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.445 5.77 0.675 ;
      RECT  0.18 1.005 4.3 1.235 ;
  END
END MDN_ND3_2
#-----------------------------------------------------------------------
#      Cell        : MDN_ND3_3
#      Description : 3-Input NAND
#      Equation    : X=!(A1&A2&A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND3_3
  CLASS CORE ;
  FOREIGN MDN_ND3_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 10.78 2.355 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 7.42 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 4.06 2.355 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 -0.14 11.37 0.14 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 1.005 11.02 1.235 ;
      RECT  7.725 1.235 7.955 3.805 ;
      RECT  1.72 3.805 11.02 4.035 ;
    END
    ANTENNADIFFAREA 9.924 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.445 10.25 0.675 ;
      RECT  1.72 1.005 7.24 1.235 ;
  END
END MDN_ND3_3
#-----------------------------------------------------------------------
#      Cell        : MDN_ND3_4
#      Description : 3-Input NAND
#      Equation    : X=!(A1&A2&A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND3_4
  CLASS CORE ;
  FOREIGN MDN_ND3_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.88 -0.14 13.61 0.14 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.405 1.005 13.26 1.235 ;
      RECT  9.405 1.235 9.635 1.565 ;
      RECT  8.845 1.565 9.635 1.795 ;
      RECT  8.845 1.795 9.075 3.805 ;
      RECT  0.18 3.805 13.26 4.035 ;
    END
    ANTENNADIFFAREA 13.232 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.445 12.49 0.675 ;
      RECT  0.18 1.005 8.78 1.235 ;
  END
END MDN_ND3_4
#-----------------------------------------------------------------------
#      Cell        : MDN_ND3_6
#      Description : 3-Input NAND
#      Equation    : X=!(A1&A2&A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND3_6
  CLASS CORE ;
  FOREIGN MDN_ND3_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 19.74 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
      RECT  18.34 2.355 18.62 2.915 ;
      RECT  19.46 2.355 19.74 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 13.02 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 6.3 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  8.4 5.46 10.195 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  19.515 -0.14 20.33 0.14 ;
      RECT  8.4 -0.14 9.52 0.14 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 0.98 19.98 1.26 ;
      RECT  13.86 1.26 14.14 1.54 ;
      RECT  13.3 1.54 14.14 1.82 ;
      RECT  13.3 1.82 13.58 3.78 ;
      RECT  0.18 3.78 19.98 4.06 ;
    END
    ANTENNADIFFAREA 19.848 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  7.67 0.445 19.21 0.675 ;
      RECT  0.18 1.005 13.26 1.235 ;
  END
END MDN_ND3_6
#-----------------------------------------------------------------------
#      Cell        : MDN_ND3_8
#      Description : 3-Input NAND
#      Equation    : X=!(A1&A2&A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND3_8
  CLASS CORE ;
  FOREIGN MDN_ND3_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 26.88 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  22.82 2.125 23.1 2.685 ;
      RECT  22.82 2.685 26.46 2.915 ;
      RECT  23.94 2.125 24.22 2.685 ;
      RECT  25.06 2.125 25.34 2.685 ;
      RECT  26.18 2.125 26.46 2.685 ;
    END
    ANTENNAGATEAREA 4.536 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.685 ;
      RECT  9.38 2.685 17.5 2.915 ;
      RECT  10.5 2.125 10.78 2.685 ;
      RECT  11.62 2.125 11.9 2.685 ;
      RECT  12.74 2.125 13.02 2.685 ;
      RECT  13.86 2.125 14.14 2.685 ;
      RECT  14.98 2.125 15.26 2.685 ;
      RECT  16.1 2.125 16.38 2.685 ;
      RECT  17.22 2.125 17.5 2.685 ;
    END
    ANTENNAGATEAREA 4.536 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 8.54 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
      RECT  2.66 2.125 2.94 2.685 ;
      RECT  3.78 2.125 4.06 2.685 ;
      RECT  4.9 2.125 5.18 2.685 ;
      RECT  6.02 2.125 6.3 2.685 ;
      RECT  7.14 2.125 7.42 2.685 ;
      RECT  8.26 2.125 8.54 2.685 ;
    END
    ANTENNAGATEAREA 4.536 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.645 5.46 27.05 5.74 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.08 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 21.84 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 16.915 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 26.88 5.74 ;
      LAYER VIA12 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  26.32 -0.14 27.05 0.14 ;
      RECT  15.12 -0.14 16.24 0.14 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 26.88 0.14 ;
      LAYER VIA12 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.31 0.935 26.645 1.305 ;
      RECT  18.31 1.305 18.65 1.535 ;
      RECT  22.215 1.305 22.585 4.295 ;
      RECT  17.735 1.535 18.65 1.875 ;
      RECT  17.735 1.875 18.11 2.1 ;
      RECT  17.735 2.1 18.105 4.295 ;
      RECT  0.18 4.295 26.7 4.665 ;
    END
    ANTENNADIFFAREA 26.464 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  9.91 0.445 25.93 0.675 ;
      RECT  0.235 0.935 17.74 1.305 ;
      RECT  18.34 2.125 18.62 2.685 ;
      RECT  18.34 2.685 21.98 2.915 ;
      RECT  19.46 2.125 19.74 2.685 ;
      RECT  20.58 2.125 20.86 2.685 ;
      RECT  21.7 2.125 21.98 2.685 ;
      RECT  21.67 5.0 23.13 5.23 ;
  END
END MDN_ND3_8
#-----------------------------------------------------------------------
#      Cell        : MDN_ND3B_1
#      Description : 3-Input NAND (A inverted input)
#      Equation    : X=!(!A&B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND3B_1
  CLASS CORE ;
  FOREIGN MDN_ND3B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 4.365 0.7 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 4.65 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  1.005 5.46 1.68 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 4.365 ;
      RECT  1.72 4.365 4.3 4.595 ;
    END
    ANTENNADIFFAREA 3.308 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.09 0.445 ;
      RECT  1.565 0.445 4.09 0.675 ;
      RECT  1.565 0.675 1.795 1.005 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  0.445 1.235 0.675 3.245 ;
      RECT  0.18 3.245 0.675 3.475 ;
      RECT  1.72 1.565 2.76 1.795 ;
  END
END MDN_ND3B_1
#-----------------------------------------------------------------------
#      Cell        : MDN_ND3B_2
#      Description : 3-Input NAND (A inverted input)
#      Equation    : X=!(!A&B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND3B_2
  CLASS CORE ;
  FOREIGN MDN_ND3B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 4.365 7.42 5.0 ;
      RECT  7.11 5.0 7.45 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.905 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 2.06 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.365 1.565 6.54 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  4.365 3.245 6.54 3.475 ;
      RECT  4.365 3.475 4.595 3.805 ;
      RECT  0.18 3.805 4.595 4.035 ;
    END
    ANTENNADIFFAREA 6.616 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 3.53 0.675 ;
      RECT  4.365 0.445 5.77 0.675 ;
      RECT  4.365 0.675 4.595 1.005 ;
      RECT  2.42 1.005 4.595 1.235 ;
      RECT  6.9 1.565 7.395 1.795 ;
      RECT  7.165 1.795 7.395 2.405 ;
      RECT  4.87 2.405 7.395 2.635 ;
      RECT  7.165 2.635 7.395 3.245 ;
      RECT  6.9 3.245 7.395 3.475 ;
  END
END MDN_ND3B_2
#-----------------------------------------------------------------------
#      Cell        : MDN_ND3B_3
#      Description : 3-Input NAND (A inverted input)
#      Equation    : X=!(!A&B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND3B_3
  CLASS CORE ;
  FOREIGN MDN_ND3B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 7.42 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 -0.14 11.37 0.14 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.44 1.005 9.075 1.235 ;
      RECT  8.845 1.235 9.075 1.565 ;
      RECT  8.845 1.565 11.02 1.795 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  8.845 3.245 11.02 3.475 ;
      RECT  8.845 3.475 9.075 4.365 ;
      RECT  0.18 4.365 9.075 4.595 ;
    END
    ANTENNADIFFAREA 9.924 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.445 10.25 0.675 ;
      RECT  0.18 1.005 7.24 1.235 ;
      RECT  3.96 1.565 8.515 1.795 ;
      RECT  8.285 1.795 8.515 2.69 ;
      RECT  4.365 1.795 4.595 3.805 ;
      RECT  3.96 3.805 4.595 4.035 ;
      RECT  9.405 2.125 10.755 2.355 ;
      RECT  9.405 2.355 9.635 2.69 ;
      RECT  10.525 2.355 10.755 2.69 ;
      RECT  8.23 5.0 9.69 5.23 ;
  END
END MDN_ND3B_3
#-----------------------------------------------------------------------
#      Cell        : MDN_ND3B_4
#      Description : 3-Input NAND (A inverted input)
#      Equation    : X=!(!A&B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND3B_4
  CLASS CORE ;
  FOREIGN MDN_ND3B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 14.14 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.765 4.365 13.26 4.595 ;
      RECT  12.765 4.595 12.995 5.46 ;
      RECT  12.765 5.46 13.44 5.74 ;
      RECT  11.38 4.365 11.875 4.595 ;
      RECT  11.645 4.595 11.875 5.46 ;
      RECT  11.2 5.46 11.875 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.765 1.005 13.26 1.235 ;
      RECT  12.765 1.235 12.995 1.565 ;
      RECT  8.845 1.565 12.995 1.795 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  8.845 3.245 12.49 3.475 ;
      RECT  8.845 3.475 9.075 4.365 ;
      RECT  0.18 4.365 9.075 4.595 ;
    END
    ANTENNADIFFAREA 12.908 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.445 12.49 0.675 ;
      RECT  0.18 1.005 8.78 1.235 ;
      RECT  13.325 1.565 13.96 1.795 ;
      RECT  13.325 1.795 13.555 2.125 ;
      RECT  9.405 2.125 13.555 2.355 ;
      RECT  9.405 2.355 9.635 2.69 ;
      RECT  10.525 2.355 10.755 2.69 ;
      RECT  11.645 2.355 11.875 2.69 ;
      RECT  12.765 2.355 12.995 2.69 ;
      RECT  13.325 2.355 13.555 3.805 ;
      RECT  13.325 3.805 13.96 4.035 ;
  END
END MDN_ND3B_4
#-----------------------------------------------------------------------
#      Cell        : MDN_ND4_1
#      Description : 4-Input NAND
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND4_1
  CLASS CORE ;
  FOREIGN MDN_ND4_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 4.65 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 1.005 4.3 1.235 ;
      RECT  3.245 1.235 3.475 4.365 ;
      RECT  0.18 4.365 4.3 4.595 ;
    END
    ANTENNADIFFAREA 4.206 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.005 2.76 1.235 ;
  END
END MDN_ND4_1
#-----------------------------------------------------------------------
#      Cell        : MDN_ND4_2
#      Description : 4-Input NAND
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND4_2
  CLASS CORE ;
  FOREIGN MDN_ND4_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.605 1.565 8.78 1.795 ;
      RECT  6.605 1.795 6.835 3.805 ;
      RECT  0.18 3.805 8.78 4.035 ;
    END
    ANTENNADIFFAREA 8.412 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.445 4.89 0.675 ;
      RECT  4.66 0.675 4.89 1.005 ;
      RECT  4.66 1.005 6.54 1.235 ;
      RECT  5.43 0.445 8.01 0.675 ;
      RECT  0.18 1.005 4.3 1.235 ;
  END
END MDN_ND4_2
#-----------------------------------------------------------------------
#      Cell        : MDN_ND4_3
#      Description : 4-Input NAND
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND4_3
  CLASS CORE ;
  FOREIGN MDN_ND4_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 13.02 2.355 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 9.66 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 6.3 2.355 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.88 -0.14 13.61 0.14 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 2.76 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 1.005 13.26 1.235 ;
      RECT  9.965 1.235 10.195 3.805 ;
      RECT  0.18 3.805 13.26 4.035 ;
    END
    ANTENNADIFFAREA 12.618 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 5.77 0.675 ;
      RECT  7.67 0.445 12.49 0.675 ;
      RECT  3.96 1.005 9.48 1.235 ;
  END
END MDN_ND4_3
#-----------------------------------------------------------------------
#      Cell        : MDN_ND4_4
#      Description : 4-Input NAND
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND4_4
  CLASS CORE ;
  FOREIGN MDN_ND4_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  17.275 -0.14 18.09 0.14 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.885 1.005 17.74 1.235 ;
      RECT  13.885 1.235 14.115 1.565 ;
      RECT  13.325 1.565 14.115 1.795 ;
      RECT  13.325 1.795 13.555 3.805 ;
      RECT  0.18 3.805 17.74 4.035 ;
    END
    ANTENNADIFFAREA 16.824 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.445 9.37 0.675 ;
      RECT  9.14 0.675 9.37 1.005 ;
      RECT  9.14 1.005 13.26 1.235 ;
      RECT  9.91 0.445 16.97 0.675 ;
      RECT  0.18 1.005 8.78 1.235 ;
  END
END MDN_ND4_4
#-----------------------------------------------------------------------
#      Cell        : MDN_ND4_6
#      Description : 4-Input NAND
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND4_6
  CLASS CORE ;
  FOREIGN MDN_ND4_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 26.88 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  20.58 2.125 26.46 2.355 ;
      RECT  20.58 2.355 20.86 2.915 ;
      RECT  21.7 2.355 21.98 2.915 ;
      RECT  22.82 2.355 23.1 2.915 ;
      RECT  23.94 2.355 24.22 2.915 ;
      RECT  25.06 2.355 25.34 2.915 ;
      RECT  26.18 2.355 26.46 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 19.74 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
      RECT  18.34 2.355 18.62 2.915 ;
      RECT  19.46 2.355 19.74 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 13.02 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 6.3 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.645 5.46 27.05 5.74 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.08 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 21.84 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 26.88 5.74 ;
      LAYER VIA12 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  26.32 -0.14 27.05 0.14 ;
      RECT  12.88 -0.14 14.0 0.14 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 26.88 0.14 ;
      LAYER VIA12 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  20.58 0.98 26.7 1.26 ;
      RECT  20.58 1.26 20.86 1.54 ;
      RECT  20.02 1.54 20.86 1.82 ;
      RECT  20.02 1.82 20.3 3.78 ;
      RECT  0.18 3.78 26.7 4.06 ;
    END
    ANTENNADIFFAREA 25.236 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  6.31 0.445 12.49 0.675 ;
      RECT  6.31 0.675 6.54 1.005 ;
      RECT  0.18 1.005 6.54 1.235 ;
      RECT  14.39 0.445 25.93 0.675 ;
      RECT  6.9 1.005 19.98 1.235 ;
  END
END MDN_ND4_6
#-----------------------------------------------------------------------
#      Cell        : MDN_ND4_8
#      Description : 4-Input NAND
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND4_8
  CLASS CORE ;
  FOREIGN MDN_ND4_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 35.84 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  27.3 2.125 35.42 2.355 ;
      RECT  27.3 2.355 27.58 2.915 ;
      RECT  28.42 2.355 28.7 2.915 ;
      RECT  29.54 2.355 29.82 2.915 ;
      RECT  30.66 2.355 30.94 2.915 ;
      RECT  31.78 2.355 32.06 2.915 ;
      RECT  32.9 2.355 33.18 2.915 ;
      RECT  34.02 2.355 34.3 2.915 ;
      RECT  35.14 2.355 35.42 2.915 ;
    END
    ANTENNAGATEAREA 4.536 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.34 2.125 18.62 2.685 ;
      RECT  18.34 2.685 26.46 2.915 ;
      RECT  19.46 2.125 19.74 2.685 ;
      RECT  20.58 2.125 20.86 2.685 ;
      RECT  21.7 2.125 21.98 2.685 ;
      RECT  22.82 2.125 23.1 2.685 ;
      RECT  23.94 2.125 24.22 2.685 ;
      RECT  25.06 2.125 25.34 2.685 ;
      RECT  26.18 2.125 26.46 2.685 ;
    END
    ANTENNAGATEAREA 4.536 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.685 ;
      RECT  9.38 2.685 17.5 2.915 ;
      RECT  10.5 2.125 10.78 2.685 ;
      RECT  11.62 2.125 11.9 2.685 ;
      RECT  12.74 2.125 13.02 2.685 ;
      RECT  13.86 2.125 14.14 2.685 ;
      RECT  14.98 2.125 15.26 2.685 ;
      RECT  16.1 2.125 16.38 2.685 ;
      RECT  17.22 2.125 17.5 2.685 ;
    END
    ANTENNAGATEAREA 4.536 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 8.54 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
      RECT  2.66 2.125 2.94 2.685 ;
      RECT  3.78 2.125 4.06 2.685 ;
      RECT  4.9 2.125 5.18 2.685 ;
      RECT  6.02 2.125 6.3 2.685 ;
      RECT  7.14 2.125 7.42 2.685 ;
      RECT  8.26 2.125 8.54 2.685 ;
    END
    ANTENNAGATEAREA 4.536 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  34.605 4.9 34.835 5.46 ;
      RECT  34.605 5.46 36.01 5.74 ;
      RECT  30.125 4.9 30.355 5.46 ;
      RECT  30.125 5.46 32.595 5.74 ;
      RECT  32.365 4.9 32.595 5.46 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.645 5.46 28.115 5.74 ;
      RECT  27.885 4.9 28.115 5.46 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 23.635 5.74 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 19.155 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 10.195 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 5.715 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 35.84 5.74 ;
      LAYER VIA12 ;
      RECT  34.87 5.47 35.13 5.73 ;
      RECT  35.43 5.47 35.69 5.73 ;
      RECT  30.39 5.47 30.65 5.73 ;
      RECT  30.95 5.47 31.21 5.73 ;
      RECT  31.51 5.47 31.77 5.73 ;
      RECT  32.07 5.47 32.33 5.73 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  27.03 5.47 27.29 5.73 ;
      RECT  27.59 5.47 27.85 5.73 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  22.55 5.47 22.81 5.73 ;
      RECT  23.11 5.47 23.37 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  18.07 5.47 18.33 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  34.72 -0.14 36.01 0.14 ;
      RECT  24.08 -0.14 25.2 0.14 ;
      RECT  15.12 -0.14 16.24 0.14 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 35.84 0.14 ;
      LAYER VIA12 ;
      RECT  34.87 -0.13 35.13 0.13 ;
      RECT  35.43 -0.13 35.69 0.13 ;
      RECT  24.23 -0.13 24.49 0.13 ;
      RECT  24.79 -0.13 25.05 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  27.255 0.935 35.66 1.305 ;
      RECT  27.255 1.305 27.625 1.495 ;
      RECT  26.695 1.495 27.625 1.865 ;
      RECT  26.695 1.865 27.065 3.735 ;
      RECT  0.18 3.735 35.66 4.105 ;
    END
    ANTENNADIFFAREA 33.648 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.55 0.445 16.97 0.675 ;
      RECT  8.55 0.675 8.78 1.005 ;
      RECT  0.18 1.005 8.78 1.235 ;
      RECT  18.87 0.445 34.89 0.675 ;
      RECT  9.14 1.005 26.7 1.235 ;
  END
END MDN_ND4_8
#-----------------------------------------------------------------------
#      Cell        : MDN_ND4B_1
#      Description : 4-Input NAND (A inverted input)
#      Equation    : X=!(!A&B1&B2&B3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND4B_1
  CLASS CORE ;
  FOREIGN MDN_ND4B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.91 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.91 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.91 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 -0.14 6.89 0.14 ;
      RECT  6.045 0.14 6.275 1.005 ;
      RECT  6.045 1.005 6.54 1.235 ;
      RECT  1.005 -0.14 1.68 0.14 ;
      RECT  1.005 0.14 1.235 0.69 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  2.685 1.235 2.915 3.805 ;
      RECT  2.42 3.805 6.54 4.035 ;
    END
    ANTENNADIFFAREA 4.206 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.565 0.37 2.97 0.6 ;
      RECT  1.565 0.6 1.795 1.565 ;
      RECT  1.565 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 3.245 ;
      RECT  1.775 3.245 2.355 3.475 ;
      RECT  1.775 3.475 2.005 4.09 ;
      RECT  3.955 1.005 5.0 1.235 ;
  END
END MDN_ND4B_1
#-----------------------------------------------------------------------
#      Cell        : MDN_ND4B_2
#      Description : 4-Input NAND (A inverted input)
#      Equation    : X=!(!A&B1&B2&B3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND4B_2
  CLASS CORE ;
  FOREIGN MDN_ND4B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 10.78 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 4.595 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  2.42 3.245 4.595 3.475 ;
      RECT  4.365 3.475 4.595 3.805 ;
      RECT  4.365 3.805 11.02 4.035 ;
    END
    ANTENNADIFFAREA 8.412 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.445 4.595 0.675 ;
      RECT  4.365 0.675 4.595 1.005 ;
      RECT  4.365 1.005 6.54 1.235 ;
      RECT  5.43 0.445 8.01 0.675 ;
      RECT  6.9 1.005 11.02 1.235 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.405 ;
      RECT  1.565 2.405 4.09 2.635 ;
      RECT  1.565 2.635 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
  END
END MDN_ND4B_2
#-----------------------------------------------------------------------
#      Cell        : MDN_ND4B_3
#      Description : 4-Input NAND (A inverted input)
#      Equation    : X=!(!A&B1&B2&B3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND4B_3
  CLASS CORE ;
  FOREIGN MDN_ND4B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.685 ;
      RECT  6.02 2.685 8.54 2.915 ;
      RECT  7.14 2.125 7.42 2.685 ;
      RECT  8.26 2.125 8.54 2.685 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 11.9 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.74 2.125 13.02 2.685 ;
      RECT  12.74 2.685 15.26 2.915 ;
      RECT  13.86 2.125 14.14 2.685 ;
      RECT  14.98 2.125 15.26 2.685 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.56 -0.14 15.85 0.14 ;
      RECT  15.005 0.14 15.235 1.005 ;
      RECT  12.92 1.005 15.5 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 3.245 ;
      RECT  2.42 3.245 5.155 3.475 ;
      RECT  4.925 3.475 5.155 3.805 ;
      RECT  4.925 3.805 15.5 4.035 ;
    END
    ANTENNADIFFAREA 12.618 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.445 8.01 0.675 ;
      RECT  9.91 0.445 14.73 0.675 ;
      RECT  6.16 1.005 11.72 1.235 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.405 ;
      RECT  1.565 2.405 4.09 2.635 ;
      RECT  1.565 2.635 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  3.75 5.0 5.21 5.23 ;
  END
END MDN_ND4B_3
#-----------------------------------------------------------------------
#      Cell        : MDN_ND4B_4
#      Description : 4-Input NAND (A inverted input)
#      Equation    : X=!(!A&B1&B2&B3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_ND4B_4
  CLASS CORE ;
  FOREIGN MDN_ND4B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 10.78 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 2.125 11.9 2.685 ;
      RECT  11.62 2.685 15.26 2.915 ;
      RECT  12.74 2.125 13.02 2.685 ;
      RECT  13.86 2.125 14.14 2.685 ;
      RECT  14.98 2.125 15.26 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  16.1 2.125 19.74 2.355 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
      RECT  18.34 2.355 18.62 2.915 ;
      RECT  19.46 2.355 19.74 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  15.12 5.46 16.915 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  11.76 5.46 12.435 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.73 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  15.12 -0.14 16.24 0.14 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 6.835 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  2.42 3.245 6.835 3.475 ;
      RECT  6.605 3.475 6.835 3.805 ;
      RECT  6.605 3.805 19.98 4.035 ;
    END
    ANTENNADIFFAREA 16.824 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.445 6.835 0.675 ;
      RECT  6.605 0.675 6.835 1.005 ;
      RECT  6.605 1.005 11.02 1.235 ;
      RECT  7.67 0.445 14.73 0.675 ;
      RECT  11.38 1.005 19.98 1.235 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.405 ;
      RECT  1.565 2.405 6.33 2.635 ;
      RECT  1.565 2.635 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
  END
END MDN_ND4B_4
#-----------------------------------------------------------------------
#      Cell        : MDN_NR2_1
#      Description : 2-Input NOR
#      Equation    : X=!(A1|A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR2_1
  CLASS CORE ;
  FOREIGN MDN_NR2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.24 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 2.24 5.74 ;
      LAYER VIA12 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.565 -0.14 2.41 0.14 ;
      RECT  1.565 0.14 1.795 1.005 ;
      RECT  1.565 1.005 2.06 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 2.24 0.14 ;
      LAYER VIA12 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 1.51 1.235 3.245 ;
      RECT  1.005 3.245 2.06 3.475 ;
    END
    ANTENNADIFFAREA 1.992 ;
  END X
END MDN_NR2_1
#-----------------------------------------------------------------------
#      Cell        : MDN_NR2_12
#      Description : 2-Input NOR
#      Equation    : X=!(A1|A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR2_12
  CLASS CORE ;
  FOREIGN MDN_NR2_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 26.88 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.95 2.125 26.46 2.355 ;
      RECT  13.95 2.355 14.37 2.38 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
      RECT  18.34 2.355 18.62 2.915 ;
      RECT  19.46 2.355 19.74 2.915 ;
      RECT  20.58 2.355 20.86 2.915 ;
      RECT  21.7 2.355 21.98 2.915 ;
      RECT  22.82 2.355 23.1 2.915 ;
      RECT  23.94 2.355 24.22 2.915 ;
      RECT  25.06 2.355 25.34 2.915 ;
      RECT  26.18 2.355 26.46 2.915 ;
      RECT  13.95 2.38 14.23 2.915 ;
    END
    ANTENNAGATEAREA 6.804 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 12.93 2.355 ;
      RECT  12.51 2.355 12.93 2.385 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.65 2.385 12.93 2.915 ;
    END
    ANTENNAGATEAREA 6.804 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  26.32 5.46 27.05 5.74 ;
      RECT  19.6 5.46 20.72 5.74 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.52 5.46 12.88 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 8.4 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 6.16 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.68 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 26.88 5.74 ;
      LAYER VIA12 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  20.31 5.47 20.57 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.2 -0.14 27.05 0.14 ;
      RECT  25.59 0.14 25.93 0.465 ;
      RECT  22.96 -0.14 24.08 0.14 ;
      RECT  23.35 0.14 23.69 0.465 ;
      RECT  20.72 -0.14 21.84 0.14 ;
      RECT  21.11 0.14 21.45 0.465 ;
      RECT  18.48 -0.14 19.6 0.14 ;
      RECT  18.87 0.14 19.21 0.465 ;
      RECT  16.24 -0.14 17.36 0.14 ;
      RECT  16.63 0.14 16.97 0.465 ;
      RECT  11.76 -0.14 15.12 0.14 ;
      RECT  12.15 0.14 12.49 0.465 ;
      RECT  14.39 0.14 14.73 0.465 ;
      RECT  9.52 -0.14 10.64 0.14 ;
      RECT  9.91 0.14 10.25 0.465 ;
      RECT  7.28 -0.14 8.4 0.14 ;
      RECT  7.67 0.14 8.01 0.465 ;
      RECT  5.04 -0.14 6.16 0.14 ;
      RECT  5.43 0.14 5.77 0.465 ;
      RECT  2.8 -0.14 3.92 0.14 ;
      RECT  3.19 0.14 3.53 0.465 ;
      RECT  -0.17 -0.14 1.68 0.14 ;
      RECT  0.95 0.14 1.29 0.465 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 26.88 0.14 ;
      LAYER VIA12 ;
      RECT  25.35 -0.13 25.61 0.13 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  23.11 -0.13 23.37 0.13 ;
      RECT  23.67 -0.13 23.93 0.13 ;
      RECT  20.87 -0.13 21.13 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 0.695 26.7 1.255 ;
      RECT  13.07 1.255 13.81 1.26 ;
      RECT  13.16 1.26 13.72 3.145 ;
      RECT  13.16 3.145 25.875 3.705 ;
    END
    ANTENNADIFFAREA 25.188 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  24.525 4.365 26.7 4.595 ;
      RECT  24.525 4.595 24.755 4.925 ;
      RECT  0.18 4.365 13.555 4.595 ;
      RECT  13.325 4.595 13.555 4.925 ;
      RECT  13.325 4.925 24.755 5.155 ;
  END
END MDN_NR2_12
#-----------------------------------------------------------------------
#      Cell        : MDN_NR2_16
#      Description : 2-Input NOR
#      Equation    : X=!(A1|A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR2_16
  CLASS CORE ;
  FOREIGN MDN_NR2_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 35.84 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.59 2.125 35.42 2.355 ;
      RECT  18.59 2.355 18.875 2.65 ;
      RECT  19.46 2.355 19.74 2.915 ;
      RECT  20.58 2.355 20.86 2.915 ;
      RECT  21.7 2.355 21.98 2.915 ;
      RECT  22.82 2.355 23.1 2.915 ;
      RECT  23.94 2.355 24.22 2.915 ;
      RECT  25.06 2.355 25.34 2.915 ;
      RECT  26.18 2.355 26.46 2.915 ;
      RECT  27.3 2.355 27.58 2.915 ;
      RECT  28.42 2.355 28.7 2.915 ;
      RECT  29.54 2.355 29.82 2.915 ;
      RECT  30.66 2.355 30.94 2.915 ;
      RECT  31.78 2.355 32.06 2.915 ;
      RECT  32.9 2.355 33.18 2.915 ;
      RECT  34.02 2.355 34.3 2.915 ;
      RECT  35.14 2.355 35.42 2.915 ;
    END
    ANTENNAGATEAREA 9.072 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 17.25 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  16.96 2.355 17.25 2.94 ;
    END
    ANTENNAGATEAREA 9.072 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  35.28 5.46 36.01 5.74 ;
      RECT  26.32 5.46 27.44 5.74 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  12.205 5.46 14.675 5.74 ;
      RECT  14.445 4.87 14.675 5.46 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 35.84 5.74 ;
      LAYER VIA12 ;
      RECT  35.43 5.47 35.69 5.73 ;
      RECT  26.47 5.47 26.73 5.73 ;
      RECT  27.03 5.47 27.29 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  13.59 5.47 13.85 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  35.16 -0.14 36.01 0.14 ;
      RECT  35.16 0.14 35.39 0.89 ;
      RECT  35.16 0.89 35.66 1.12 ;
      RECT  33.6 -0.14 34.275 0.14 ;
      RECT  34.045 0.14 34.275 0.89 ;
      RECT  33.78 0.89 34.275 1.12 ;
      RECT  31.92 -0.14 32.595 0.14 ;
      RECT  32.365 0.14 32.595 0.52 ;
      RECT  30.125 -0.14 30.8 0.14 ;
      RECT  30.125 0.14 30.355 0.52 ;
      RECT  25.645 -0.14 28.115 0.14 ;
      RECT  25.645 0.14 25.875 0.52 ;
      RECT  27.885 0.14 28.115 0.52 ;
      RECT  22.96 -0.14 23.635 0.14 ;
      RECT  23.405 0.14 23.635 0.52 ;
      RECT  21.165 -0.14 21.84 0.14 ;
      RECT  21.165 0.14 21.395 0.52 ;
      RECT  18.48 -0.14 19.155 0.14 ;
      RECT  18.925 0.14 19.155 0.52 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.52 ;
      RECT  12.205 -0.14 14.675 0.14 ;
      RECT  12.205 0.14 12.435 0.52 ;
      RECT  14.445 0.14 14.675 0.52 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.52 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.52 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.52 ;
      RECT  1.565 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.52 ;
      RECT  1.565 0.14 1.795 0.89 ;
      RECT  1.565 0.89 2.06 1.12 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 0.89 ;
      RECT  0.18 0.89 0.675 1.12 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 35.84 0.14 ;
      LAYER VIA12 ;
      RECT  35.43 -0.13 35.69 0.13 ;
      RECT  33.75 -0.13 34.01 0.13 ;
      RECT  32.07 -0.13 32.33 0.13 ;
      RECT  30.39 -0.13 30.65 0.13 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  27.03 -0.13 27.29 0.13 ;
      RECT  27.59 -0.13 27.85 0.13 ;
      RECT  23.11 -0.13 23.37 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  18.63 -0.13 18.89 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  13.59 -0.13 13.85 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 33.42 1.35 ;
      RECT  1.005 1.35 34.835 1.745 ;
      RECT  1.005 1.745 3.17 1.87 ;
      RECT  32.67 1.745 34.835 1.87 ;
      RECT  17.55 1.745 18.29 3.245 ;
      RECT  17.55 3.245 34.835 3.985 ;
    END
    ANTENNADIFFAREA 33.424 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  33.485 4.365 35.66 4.595 ;
      RECT  33.485 4.595 33.715 4.925 ;
      RECT  0.18 4.365 18.035 4.595 ;
      RECT  17.805 4.595 18.035 4.925 ;
      RECT  17.805 4.925 33.715 5.155 ;
  END
END MDN_NR2_16
#-----------------------------------------------------------------------
#      Cell        : MDN_NR2_2
#      Description : 2-Input NOR
#      Equation    : X=!(A1|A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR2_2
  CLASS CORE ;
  FOREIGN MDN_NR2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.685 ;
      RECT  2.66 2.685 4.06 2.915 ;
      RECT  3.78 2.125 4.06 2.685 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 1.82 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 4.65 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  2.125 1.235 2.355 3.245 ;
      RECT  2.125 3.245 3.53 3.475 ;
    END
    ANTENNADIFFAREA 3.928 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  2.42 4.365 4.3 4.595 ;
      RECT  2.685 4.595 2.915 4.925 ;
      RECT  0.95 4.925 2.915 5.155 ;
  END
END MDN_NR2_2
#-----------------------------------------------------------------------
#      Cell        : MDN_NR2_3
#      Description : 2-Input NOR
#      Equation    : X=!(A1|A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR2_3
  CLASS CORE ;
  FOREIGN MDN_NR2_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 6.3 2.355 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 6.54 1.235 ;
      RECT  3.245 1.235 3.475 4.365 ;
      RECT  3.245 4.365 6.54 4.595 ;
    END
    ANTENNADIFFAREA 6.378 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 4.925 5.77 5.155 ;
  END
END MDN_NR2_3
#-----------------------------------------------------------------------
#      Cell        : MDN_NR2_4
#      Description : 2-Input NOR
#      Equation    : X=!(A1|A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR2_4
  CLASS CORE ;
  FOREIGN MDN_NR2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.685 ;
      RECT  4.9 2.685 8.54 2.915 ;
      RECT  6.02 2.125 6.3 2.685 ;
      RECT  7.14 2.125 7.42 2.685 ;
      RECT  8.26 2.125 8.54 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 4.06 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
      RECT  2.66 2.125 2.94 2.685 ;
      RECT  3.78 2.125 4.06 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 3.475 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 8.78 1.235 ;
      RECT  4.365 1.235 4.595 3.245 ;
      RECT  4.365 3.245 8.01 3.475 ;
    END
    ANTENNADIFFAREA 8.18 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  6.605 4.365 8.78 4.595 ;
      RECT  6.605 4.595 6.835 4.925 ;
      RECT  0.18 4.365 4.595 4.595 ;
      RECT  4.365 4.595 4.595 4.925 ;
      RECT  4.365 4.925 6.835 5.155 ;
  END
END MDN_NR2_4
#-----------------------------------------------------------------------
#      Cell        : MDN_NR2_6
#      Description : 2-Input NOR
#      Equation    : X=!(A1|A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR2_6
  CLASS CORE ;
  FOREIGN MDN_NR2_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 7.42 2.685 ;
      RECT  7.14 2.685 13.02 2.915 ;
      RECT  8.26 2.125 8.54 2.685 ;
      RECT  9.38 2.125 9.66 2.685 ;
      RECT  10.5 2.125 10.78 2.685 ;
      RECT  11.62 2.125 11.9 2.685 ;
      RECT  12.74 2.125 13.02 2.685 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 6.3 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.88 5.46 13.61 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 0.98 13.26 1.26 ;
      RECT  6.58 1.26 6.86 3.78 ;
      RECT  6.58 3.78 12.49 4.06 ;
    END
    ANTENNADIFFAREA 12.432 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  11.085 4.365 13.26 4.595 ;
      RECT  11.085 4.595 11.315 4.925 ;
      RECT  0.18 4.365 6.835 4.595 ;
      RECT  6.605 4.595 6.835 4.925 ;
      RECT  6.605 4.925 11.315 5.155 ;
  END
END MDN_NR2_6
#-----------------------------------------------------------------------
#      Cell        : MDN_NR2_8
#      Description : 2-Input NOR
#      Equation    : X=!(A1|A2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR2_8
  CLASS CORE ;
  FOREIGN MDN_NR2_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.685 ;
      RECT  9.38 2.685 17.5 2.915 ;
      RECT  10.5 2.125 10.78 2.685 ;
      RECT  11.62 2.125 11.9 2.685 ;
      RECT  12.74 2.125 13.02 2.685 ;
      RECT  13.86 2.125 14.14 2.685 ;
      RECT  14.98 2.125 15.26 2.685 ;
      RECT  16.1 2.125 16.38 2.685 ;
      RECT  17.22 2.125 17.5 2.685 ;
    END
    ANTENNAGATEAREA 4.536 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 8.54 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 4.536 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  17.36 5.46 18.09 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.635 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.635 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.635 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.635 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.635 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.635 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.635 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.635 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 0.865 17.74 1.235 ;
      RECT  8.59 1.235 9.33 1.26 ;
      RECT  8.775 1.26 9.145 3.75 ;
      RECT  8.775 3.75 9.35 4.09 ;
      RECT  9.01 4.09 9.35 4.295 ;
      RECT  9.01 4.295 17.685 4.665 ;
    END
    ANTENNADIFFAREA 17.008 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 4.365 8.78 4.595 ;
      RECT  8.55 4.595 8.78 4.925 ;
      RECT  8.55 4.925 16.97 5.155 ;
  END
END MDN_NR2_8
#-----------------------------------------------------------------------
#      Cell        : MDN_NR2B_1
#      Description : 2-Input NOR (A inverted input)
#      Equation    : X=!(!A|B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR2B_1
  CLASS CORE ;
  FOREIGN MDN_NR2B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 4.65 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  0.56 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 4.3 1.235 ;
      RECT  2.685 1.235 2.915 3.805 ;
      RECT  2.42 3.805 2.915 4.035 ;
    END
    ANTENNADIFFAREA 2.126 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  2.63 0.37 2.97 0.445 ;
      RECT  1.565 0.445 2.97 0.675 ;
      RECT  1.565 0.675 1.795 1.565 ;
      RECT  1.565 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 3.245 ;
      RECT  1.72 3.245 2.355 3.475 ;
  END
END MDN_NR2B_1
#-----------------------------------------------------------------------
#      Cell        : MDN_NR2B_2
#      Description : 2-Input NOR (A inverted input)
#      Equation    : X=!(!A|B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR2B_2
  CLASS CORE ;
  FOREIGN MDN_NR2B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 4.365 6.54 4.595 ;
      RECT  6.045 4.595 6.275 5.46 ;
      RECT  5.6 5.46 6.89 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 6.89 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 6.54 1.235 ;
      RECT  4.365 1.235 4.595 3.245 ;
      RECT  3.19 3.245 4.595 3.475 ;
    END
    ANTENNADIFFAREA 3.928 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 2.405 ;
      RECT  2.125 2.405 4.09 2.635 ;
      RECT  2.125 2.635 2.355 3.245 ;
      RECT  1.72 3.245 2.355 3.475 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 4.925 ;
      RECT  2.42 4.365 2.915 4.595 ;
      RECT  2.685 4.595 2.915 4.925 ;
      RECT  2.685 4.925 5.77 5.155 ;
  END
END MDN_NR2B_2
#-----------------------------------------------------------------------
#      Cell        : MDN_NR2B_3
#      Description : 2-Input NOR (A inverted input)
#      Equation    : X=!(!A|B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR2B_3
  CLASS CORE ;
  FOREIGN MDN_NR2B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 8.54 2.355 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 4.365 8.78 4.595 ;
      RECT  8.285 4.595 8.515 5.46 ;
      RECT  7.84 5.46 9.13 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 8.78 1.235 ;
      RECT  5.485 1.235 5.715 3.245 ;
      RECT  3.19 3.245 5.715 3.475 ;
    END
    ANTENNADIFFAREA 6.054 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 2.685 ;
      RECT  2.125 2.685 5.155 2.915 ;
      RECT  2.685 2.35 2.915 2.685 ;
      RECT  3.805 2.35 4.035 2.685 ;
      RECT  4.925 2.35 5.155 2.685 ;
      RECT  2.125 2.915 2.355 3.245 ;
      RECT  1.72 3.245 2.355 3.475 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 4.925 ;
      RECT  2.42 4.365 2.915 4.595 ;
      RECT  2.685 4.595 2.915 4.925 ;
      RECT  2.685 4.925 8.01 5.155 ;
  END
END MDN_NR2B_3
#-----------------------------------------------------------------------
#      Cell        : MDN_NR2B_4
#      Description : 2-Input NOR (A inverted input)
#      Equation    : X=!(!A|B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR2B_4
  CLASS CORE ;
  FOREIGN MDN_NR2B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 10.78 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 11.02 1.235 ;
      RECT  6.605 1.235 6.835 3.245 ;
      RECT  3.19 3.245 6.835 3.475 ;
    END
    ANTENNADIFFAREA 8.18 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 2.405 ;
      RECT  2.125 2.405 6.33 2.635 ;
      RECT  2.125 2.635 2.355 3.245 ;
      RECT  1.72 3.245 2.355 3.475 ;
      RECT  6.605 4.365 11.02 4.595 ;
      RECT  6.605 4.595 6.835 4.925 ;
      RECT  2.42 4.365 4.595 4.595 ;
      RECT  4.365 4.595 4.595 4.925 ;
      RECT  4.365 4.925 6.835 5.155 ;
  END
END MDN_NR2B_4
#-----------------------------------------------------------------------
#      Cell        : MDN_NR3_1
#      Description : 3-Input NOR
#      Equation    : X=!(A1|A2|A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR3_1
  CLASS CORE ;
  FOREIGN MDN_NR3_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      RECT  3.245 0.14 3.475 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 3.53 ;
    END
    ANTENNADIFFAREA 3.314 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 4.365 2.76 4.595 ;
  END
END MDN_NR3_1
#-----------------------------------------------------------------------
#      Cell        : MDN_NR3_2
#      Description : 3-Input NOR
#      Equation    : X=!(A1|A2|A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR3_2
  CLASS CORE ;
  FOREIGN MDN_NR3_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 6.54 1.235 ;
      RECT  4.365 1.235 4.595 3.245 ;
      RECT  4.365 3.245 5.77 3.475 ;
    END
    ANTENNADIFFAREA 5.156 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  1.83 4.595 2.06 4.925 ;
      RECT  1.83 4.925 3.53 5.155 ;
      RECT  6.045 4.365 6.54 4.595 ;
      RECT  6.045 4.595 6.275 4.925 ;
      RECT  2.42 4.365 5.155 4.595 ;
      RECT  4.925 4.595 5.155 4.925 ;
      RECT  4.925 4.925 6.275 5.155 ;
  END
END MDN_NR3_2
#-----------------------------------------------------------------------
#      Cell        : MDN_NR3_3
#      Description : 3-Input NOR
#      Equation    : X=!(A1|A2|A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR3_3
  CLASS CORE ;
  FOREIGN MDN_NR3_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 10.78 2.355 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 7.42 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 4.06 2.355 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 5.46 11.37 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.72 1.005 11.02 1.235 ;
      RECT  7.725 1.235 7.955 3.245 ;
      RECT  7.725 3.245 10.25 3.475 ;
    END
    ANTENNADIFFAREA 7.896 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 4.365 7.24 4.595 ;
      RECT  10.525 4.365 11.02 4.595 ;
      RECT  10.525 4.595 10.755 4.925 ;
      RECT  9.14 4.365 9.635 4.595 ;
      RECT  9.405 4.595 9.635 4.925 ;
      RECT  5.43 4.925 10.755 5.155 ;
  END
END MDN_NR3_3
#-----------------------------------------------------------------------
#      Cell        : MDN_NR3_4
#      Description : 3-Input NOR
#      Equation    : X=!(A1|A2|A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR3_4
  CLASS CORE ;
  FOREIGN MDN_NR3_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.88 5.46 13.61 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 13.26 1.235 ;
      RECT  8.845 1.235 9.075 3.245 ;
      RECT  8.845 3.245 12.49 3.475 ;
    END
    ANTENNADIFFAREA 10.636 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 4.365 8.78 4.595 ;
      RECT  12.765 4.365 13.26 4.595 ;
      RECT  12.765 4.595 12.995 4.925 ;
      RECT  11.38 4.365 11.875 4.595 ;
      RECT  11.645 4.595 11.875 4.925 ;
      RECT  5.43 4.925 12.995 5.155 ;
  END
END MDN_NR3_4
#-----------------------------------------------------------------------
#      Cell        : MDN_NR3_6
#      Description : 3-Input NOR
#      Equation    : X=!(A1|A2|A3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR3_6
  CLASS CORE ;
  FOREIGN MDN_NR3_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 19.74 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
      RECT  18.34 2.355 18.62 2.915 ;
      RECT  19.46 2.355 19.74 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 13.02 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 6.3 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 3.402 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  19.6 5.46 20.33 5.74 ;
      RECT  8.4 5.46 9.52 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  11.76 -0.14 12.435 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  7.725 -0.14 10.195 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 0.98 19.98 1.26 ;
      RECT  13.3 1.26 13.58 3.22 ;
      RECT  13.3 3.22 19.21 3.5 ;
    END
    ANTENNADIFFAREA 16.116 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 4.365 13.26 4.595 ;
      RECT  19.485 4.365 19.98 4.595 ;
      RECT  19.485 4.595 19.715 4.925 ;
      RECT  18.1 4.365 18.6 4.595 ;
      RECT  18.37 4.595 18.6 4.925 ;
      RECT  7.67 4.925 19.715 5.155 ;
  END
END MDN_NR3_6
#-----------------------------------------------------------------------
#      Cell        : MDN_NR3B_1
#      Description : 3-Input NOR (A inverted input)
#      Equation    : X=!(!A|B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR3B_1
  CLASS CORE ;
  FOREIGN MDN_NR3B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.72 1.005 4.3 1.235 ;
      RECT  3.805 1.235 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
    END
    ANTENNADIFFAREA 2.74 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 1.795 4.595 ;
      RECT  1.565 4.595 1.795 4.925 ;
      RECT  1.565 4.925 4.09 5.155 ;
      RECT  3.75 5.155 4.09 5.23 ;
      RECT  1.72 3.805 2.355 4.035 ;
      RECT  2.125 4.035 2.355 4.365 ;
      RECT  2.125 4.365 2.76 4.595 ;
  END
END MDN_NR3B_1
#-----------------------------------------------------------------------
#      Cell        : MDN_NR3B_2
#      Description : 3-Input NOR (A inverted input)
#      Equation    : X=!(!A|B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR3B_2
  CLASS CORE ;
  FOREIGN MDN_NR3B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 4.365 7.42 5.0 ;
      RECT  7.11 5.0 7.45 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 9.13 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 4.595 1.235 ;
      RECT  4.365 1.235 4.595 1.565 ;
      RECT  4.365 1.565 6.54 1.795 ;
      RECT  5.485 1.795 5.715 3.53 ;
    END
    ANTENNADIFFAREA 5.156 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  4.98 1.005 7.395 1.235 ;
      RECT  7.165 1.235 7.395 3.245 ;
      RECT  6.9 3.245 7.395 3.475 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  6.045 4.365 6.54 4.595 ;
      RECT  6.045 4.595 6.275 4.925 ;
      RECT  4.66 4.365 5.155 4.595 ;
      RECT  4.925 4.595 5.155 4.925 ;
      RECT  3.19 4.925 6.275 5.155 ;
  END
END MDN_NR3B_2
#-----------------------------------------------------------------------
#      Cell        : MDN_NR3B_3
#      Description : 3-Input NOR (A inverted input)
#      Equation    : X=!(!A|B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR3B_3
  CLASS CORE ;
  FOREIGN MDN_NR3B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 7.42 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 5.46 11.37 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 9.075 1.235 ;
      RECT  8.845 1.235 9.075 1.565 ;
      RECT  8.845 1.565 11.02 1.795 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  8.44 3.245 11.02 3.475 ;
    END
    ANTENNADIFFAREA 8.22 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 9.69 0.6 ;
      RECT  3.96 1.565 8.515 1.795 ;
      RECT  8.285 1.795 8.515 2.69 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  3.96 3.245 4.595 3.475 ;
      RECT  9.515 2.405 10.81 2.635 ;
      RECT  0.18 4.365 7.24 4.595 ;
      RECT  5.43 4.925 10.25 5.155 ;
  END
END MDN_NR3B_3
#-----------------------------------------------------------------------
#      Cell        : MDN_NR3B_4
#      Description : 3-Input NOR (A inverted input)
#      Equation    : X=!(!A|B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR3B_4
  CLASS CORE ;
  FOREIGN MDN_NR3B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 4.365 14.14 5.0 ;
      RECT  13.83 5.0 14.17 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 11.315 1.235 ;
      RECT  11.085 1.235 11.315 1.565 ;
      RECT  11.085 1.565 13.26 1.795 ;
      RECT  11.085 1.795 11.315 3.245 ;
      RECT  9.14 3.245 13.26 3.475 ;
    END
    ANTENNADIFFAREA 10.96 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 11.93 0.6 ;
      RECT  13.62 1.565 14.115 1.795 ;
      RECT  13.885 1.795 14.115 2.405 ;
      RECT  11.59 2.405 14.115 2.635 ;
      RECT  13.885 2.635 14.115 3.245 ;
      RECT  13.62 3.245 14.115 3.475 ;
      RECT  9.35 2.405 10.81 2.635 ;
      RECT  0.18 4.365 8.78 4.595 ;
      RECT  5.43 4.925 12.49 5.155 ;
  END
END MDN_NR3B_4
#-----------------------------------------------------------------------
#      Cell        : MDN_NR4_1
#      Description : 4-Input NOR
#      Equation    : X=!(A1|A2|A3|A4)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR4_1
  CLASS CORE ;
  FOREIGN MDN_NR4_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 4.65 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  3.245 1.235 3.475 4.365 ;
      RECT  3.245 4.365 4.3 4.595 ;
    END
    ANTENNADIFFAREA 3.354 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 4.365 2.76 4.595 ;
  END
END MDN_NR4_1
#-----------------------------------------------------------------------
#      Cell        : MDN_NR4_2
#      Description : 4-Input NOR
#      Equation    : X=!(A1|A2|A3|A4)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR4_2
  CLASS CORE ;
  FOREIGN MDN_NR4_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      RECT  3.245 0.14 3.475 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 8.78 1.235 ;
      RECT  6.605 1.235 6.835 3.245 ;
      RECT  6.605 3.245 8.01 3.475 ;
    END
    ANTENNADIFFAREA 6.384 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  2.42 4.365 6.54 4.595 ;
      RECT  8.285 4.365 8.78 4.595 ;
      RECT  8.285 4.595 8.515 4.925 ;
      RECT  6.9 4.365 7.395 4.595 ;
      RECT  7.165 4.595 7.395 4.925 ;
      RECT  5.43 4.925 8.515 5.155 ;
      RECT  0.95 4.925 3.53 5.155 ;
  END
END MDN_NR4_2
#-----------------------------------------------------------------------
#      Cell        : MDN_NR4_3
#      Description : 4-Input NOR
#      Equation    : X=!(A1|A2|A3|A4)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR4_3
  CLASS CORE ;
  FOREIGN MDN_NR4_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.685 ;
      RECT  10.5 2.685 13.02 2.915 ;
      RECT  11.62 2.125 11.9 2.685 ;
      RECT  12.74 2.125 13.02 2.685 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 9.66 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.685 ;
      RECT  3.78 2.685 6.3 2.915 ;
      RECT  4.9 2.125 5.18 2.685 ;
      RECT  6.02 2.125 6.3 2.685 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.88 5.46 13.61 5.74 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 13.26 1.235 ;
      RECT  9.965 1.235 10.195 3.805 ;
      RECT  9.965 3.805 12.49 4.035 ;
    END
    ANTENNADIFFAREA 9.738 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.96 4.365 9.48 4.595 ;
      RECT  12.765 4.365 13.26 4.595 ;
      RECT  12.765 4.595 12.995 4.925 ;
      RECT  11.38 4.365 11.875 4.595 ;
      RECT  11.645 4.595 11.875 4.925 ;
      RECT  7.67 4.925 12.995 5.155 ;
      RECT  0.95 4.925 5.77 5.155 ;
  END
END MDN_NR4_3
#-----------------------------------------------------------------------
#      Cell        : MDN_NR4_4
#      Description : 4-Input NOR
#      Equation    : X=!(A1|A2|A3|A4)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR4_4
  CLASS CORE ;
  FOREIGN MDN_NR4_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
      RECT  13.86 2.355 14.14 2.92 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  17.36 5.46 18.09 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.14 1.005 17.74 1.235 ;
      RECT  13.325 1.235 13.555 3.245 ;
      RECT  13.325 3.245 16.97 3.475 ;
    END
    ANTENNADIFFAREA 13.092 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 4.365 8.78 4.595 ;
      RECT  17.245 4.365 17.74 4.595 ;
      RECT  17.245 4.595 17.475 4.925 ;
      RECT  15.86 4.365 16.355 4.595 ;
      RECT  16.125 4.595 16.355 4.925 ;
      RECT  9.1 4.365 13.555 4.595 ;
      RECT  13.325 4.595 13.555 4.925 ;
      RECT  13.325 4.925 17.475 5.155 ;
      RECT  5.43 4.925 12.49 5.155 ;
  END
END MDN_NR4_4
#-----------------------------------------------------------------------
#      Cell        : MDN_NR4B_1
#      Description : 4-Input NOR (A inverted input)
#      Equation    : X=!(!A|B1|B2|B3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR4B_1
  CLASS CORE ;
  FOREIGN MDN_NR4B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 4.365 5.18 5.0 ;
      RECT  4.87 5.0 5.21 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  3.805 1.235 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
    END
    ANTENNADIFFAREA 3.354 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.09 0.445 ;
      RECT  3.75 0.445 4.85 0.675 ;
      RECT  4.62 0.675 4.85 1.005 ;
      RECT  4.62 1.005 5.155 1.235 ;
      RECT  4.925 1.235 5.155 3.245 ;
      RECT  4.66 3.245 5.155 3.475 ;
      RECT  1.72 4.365 2.76 4.595 ;
  END
END MDN_NR4B_1
#-----------------------------------------------------------------------
#      Cell        : MDN_NR4B_2
#      Description : 4-Input NOR (A inverted input)
#      Equation    : X=!(!A|B1|B2|B3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR4B_2
  CLASS CORE ;
  FOREIGN MDN_NR4B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 4.365 9.66 5.0 ;
      RECT  9.35 5.0 9.69 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 6.835 1.235 ;
      RECT  6.605 1.235 6.835 1.565 ;
      RECT  6.605 1.565 8.78 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  6.605 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 6.708 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  9.14 1.565 9.635 1.795 ;
      RECT  9.405 1.795 9.635 2.405 ;
      RECT  7.11 2.405 9.635 2.635 ;
      RECT  9.405 2.635 9.635 3.245 ;
      RECT  9.14 3.245 9.635 3.475 ;
      RECT  2.42 4.365 6.54 4.595 ;
      RECT  0.95 4.925 3.53 5.155 ;
      RECT  5.43 4.925 8.01 5.155 ;
  END
END MDN_NR4B_2
#-----------------------------------------------------------------------
#      Cell        : MDN_NR4B_3
#      Description : 4-Input NOR (A inverted input)
#      Equation    : X=!(!A|B1|B2|B3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR4B_3
  CLASS CORE ;
  FOREIGN MDN_NR4B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 4.365 14.14 5.0 ;
      RECT  13.83 5.0 14.17 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 9.66 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 6.3 2.355 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  11.76 -0.14 12.435 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 10.195 1.235 ;
      RECT  9.965 1.235 10.195 1.565 ;
      RECT  9.965 1.565 13.26 1.795 ;
      RECT  9.965 1.795 10.195 3.245 ;
      RECT  9.965 3.245 13.26 3.475 ;
    END
    ANTENNADIFFAREA 10.062 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  13.62 1.565 14.115 1.795 ;
      RECT  13.885 1.795 14.115 2.405 ;
      RECT  10.47 2.405 14.115 2.635 ;
      RECT  13.885 2.635 14.115 3.245 ;
      RECT  13.62 3.245 14.115 3.475 ;
      RECT  3.96 4.365 9.48 4.595 ;
      RECT  0.95 4.925 5.77 5.155 ;
      RECT  7.67 4.925 12.49 5.155 ;
  END
END MDN_NR4B_3
#-----------------------------------------------------------------------
#      Cell        : MDN_NR4B_4
#      Description : 4-Input NOR (A inverted input)
#      Equation    : X=!(!A|B1|B2|B3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_NR4B_4
  CLASS CORE ;
  FOREIGN MDN_NR4B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.34 4.365 18.62 5.0 ;
      RECT  18.31 5.0 18.65 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  8.4 5.46 9.52 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  7.725 -0.14 10.195 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 13.555 1.235 ;
      RECT  13.325 1.235 13.555 1.565 ;
      RECT  13.325 1.565 17.74 1.795 ;
      RECT  13.325 1.795 13.555 3.245 ;
      RECT  13.325 3.245 17.74 3.475 ;
    END
    ANTENNADIFFAREA 13.416 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  18.1 1.565 18.595 1.795 ;
      RECT  18.365 1.795 18.595 2.405 ;
      RECT  13.83 2.405 18.595 2.635 ;
      RECT  18.365 2.635 18.595 3.245 ;
      RECT  18.1 3.245 18.595 3.475 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.07 4.595 4.3 4.925 ;
      RECT  4.07 4.925 8.01 5.155 ;
      RECT  4.66 4.365 13.26 4.595 ;
      RECT  9.91 4.925 16.97 5.155 ;
  END
END MDN_NR4B_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OA2111_1
#      Description : One 2-input OR into 4-input AND
#      Equation    : X=(A1|A2)&B1&B2&B3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA2111_1
  CLASS CORE ;
  FOREIGN MDN_OA2111_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 6.89 0.14 ;
      RECT  5.485 0.14 5.715 1.565 ;
      RECT  3.96 1.565 5.715 1.795 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.19 1.005 5.0 1.235 ;
      RECT  4.365 3.805 5.0 4.035 ;
      RECT  4.365 4.035 4.595 4.365 ;
      RECT  3.96 4.365 4.595 4.595 ;
      RECT  4.925 4.365 6.22 4.595 ;
      RECT  4.925 4.595 5.155 4.925 ;
      RECT  5.99 4.595 6.22 5.0 ;
      RECT  1.72 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 4.925 ;
      RECT  0.95 4.925 5.155 5.155 ;
      RECT  5.99 5.0 6.33 5.23 ;
  END
END MDN_OA2111_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OA2111_2
#      Description : One 2-input OR into 4-input AND
#      Equation    : X=(A1|A2)&B1&B2&B3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA2111_2
  CLASS CORE ;
  FOREIGN MDN_OA2111_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  8.4 5.46 9.13 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 1.565 ;
      RECT  3.96 1.565 5.715 1.795 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  6.2 3.245 7.24 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.19 0.445 4.595 0.675 ;
      RECT  4.365 0.675 4.595 1.005 ;
      RECT  4.365 1.005 5.0 1.235 ;
      RECT  1.72 1.565 2.76 1.795 ;
      RECT  4.365 3.805 5.0 4.035 ;
      RECT  4.365 4.035 4.595 4.365 ;
      RECT  3.96 4.365 4.595 4.595 ;
      RECT  4.925 4.365 6.22 4.595 ;
      RECT  4.925 4.595 5.155 4.925 ;
      RECT  5.99 4.595 6.22 5.0 ;
      RECT  0.18 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 4.925 ;
      RECT  0.95 4.925 5.155 5.155 ;
      RECT  5.99 5.0 7.45 5.23 ;
  END
END MDN_OA2111_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OA2111_4
#      Description : One 2-input OR into 4-input AND
#      Equation    : X=(A1|A2)&B1&B2&B3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA2111_4
  CLASS CORE ;
  FOREIGN MDN_OA2111_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 1.565 ;
      RECT  3.96 1.565 5.715 1.795 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 10.195 1.795 ;
      RECT  9.965 1.795 10.195 3.245 ;
      RECT  6.2 3.245 10.195 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.19 1.005 5.0 1.235 ;
      RECT  7.165 2.35 7.395 2.685 ;
      RECT  7.165 2.685 9.635 2.915 ;
      RECT  8.285 2.35 8.515 2.685 ;
      RECT  9.405 2.35 9.635 2.685 ;
      RECT  4.365 3.805 5.0 4.035 ;
      RECT  4.365 4.035 4.595 4.365 ;
      RECT  3.96 4.365 4.595 4.595 ;
      RECT  4.925 4.365 6.22 4.595 ;
      RECT  4.925 4.595 5.155 4.925 ;
      RECT  5.99 4.595 6.22 5.0 ;
      RECT  1.72 1.565 3.475 1.795 ;
      RECT  3.245 1.795 3.475 4.925 ;
      RECT  0.95 4.925 5.155 5.155 ;
      RECT  5.99 5.0 7.45 5.23 ;
  END
END MDN_OA2111_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OA211_1
#      Description : One 2-input OR into 3-input AND
#      Equation    : X=(A1|A2)&B1&B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA211_1
  CLASS CORE ;
  FOREIGN MDN_OA211_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.005 5.715 1.235 ;
      RECT  5.485 1.235 5.715 3.805 ;
      RECT  4.66 3.805 5.715 4.035 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 3.245 ;
      RECT  3.805 3.245 5.155 3.475 ;
      RECT  3.805 3.475 4.035 3.805 ;
      RECT  1.72 3.805 4.035 4.035 ;
  END
END MDN_OA211_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OA211_2
#      Description : One 2-input OR into 3-input AND
#      Equation    : X=(A1|A2)&B1&B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA211_2
  CLASS CORE ;
  FOREIGN MDN_OA211_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.75 0.37 4.09 0.6 ;
      RECT  3.78 0.6 4.06 1.235 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 6.54 1.795 ;
      RECT  5.485 1.795 5.715 3.805 ;
      RECT  4.66 3.805 6.54 4.035 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  4.98 1.005 6.22 1.235 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.805 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 2.405 ;
      RECT  3.805 2.405 5.21 2.635 ;
      RECT  3.805 2.635 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
      RECT  3.805 3.475 4.035 3.805 ;
      RECT  1.72 3.805 4.035 4.035 ;
  END
END MDN_OA211_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OA211_4
#      Description : One 2-input OR into 3-input AND
#      Equation    : X=(A1|A2)&B1&B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA211_4
  CLASS CORE ;
  FOREIGN MDN_OA211_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.005 5.715 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  5.485 1.565 8.78 1.795 ;
      RECT  6.605 1.795 6.835 3.805 ;
      RECT  4.66 3.805 8.78 4.035 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  0.18 1.005 2.76 1.235 ;
      RECT  3.96 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 2.405 ;
      RECT  4.925 2.405 6.33 2.635 ;
      RECT  4.925 2.635 5.155 3.25 ;
      RECT  3.96 3.245 4.3 3.25 ;
      RECT  3.805 3.25 5.155 3.48 ;
      RECT  3.805 3.48 4.035 3.805 ;
      RECT  1.72 3.805 4.035 4.035 ;
      RECT  7.165 2.35 7.395 2.685 ;
      RECT  7.165 2.685 8.515 2.915 ;
      RECT  8.285 2.35 8.515 2.685 ;
  END
END MDN_OA211_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OA21_1
#      Description : One 2-input OR into 2-input AND
#      Equation    : X=(A1|A2)&B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA21_1
  CLASS CORE ;
  FOREIGN MDN_OA21_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.445 1.005 2.06 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.09 0.6 ;
      RECT  3.75 0.6 3.98 1.005 ;
      RECT  3.245 1.005 3.98 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  0.18 1.565 3.475 1.795 ;
      RECT  1.005 1.795 1.235 3.5 ;
      RECT  0.95 0.445 2.705 0.675 ;
      RECT  2.475 0.675 2.705 1.29 ;
      RECT  1.72 4.365 2.76 4.595 ;
  END
END MDN_OA21_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OA21_2
#      Description : One 2-input OR into 2-input AND
#      Equation    : X=(A1|A2)&B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA21_2
  CLASS CORE ;
  FOREIGN MDN_OA21_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.445 1.005 2.06 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.96 1.565 5.0 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  3.96 3.245 5.0 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  3.75 0.6 3.98 1.005 ;
      RECT  3.245 1.005 3.98 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  0.18 1.565 3.475 1.795 ;
      RECT  1.005 1.795 1.235 3.53 ;
      RECT  0.95 0.445 2.705 0.675 ;
      RECT  2.475 0.675 2.705 1.29 ;
      RECT  1.72 4.365 2.76 4.595 ;
  END
END MDN_OA21_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OA21_3
#      Description : One 2-input OR into 2-input AND
#      Equation    : X=(A1|A2)&B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA21_3
  CLASS CORE ;
  FOREIGN MDN_OA21_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.18 4.365 0.66 4.595 ;
      RECT  0.43 4.595 0.66 5.46 ;
      RECT  -0.17 5.46 0.66 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 6.89 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.445 1.005 2.06 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.96 1.565 6.54 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  3.96 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 4.536 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  3.75 0.6 3.98 1.005 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  3.245 1.005 3.98 1.235 ;
      RECT  4.98 1.005 6.22 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  0.18 1.565 3.475 1.795 ;
      RECT  1.005 1.795 1.235 3.5 ;
      RECT  0.95 0.445 2.705 0.675 ;
      RECT  2.475 0.675 2.705 1.29 ;
      RECT  1.72 4.365 2.76 4.595 ;
  END
END MDN_OA21_3
#-----------------------------------------------------------------------
#      Cell        : MDN_OA21_4
#      Description : One 2-input OR into 2-input AND
#      Equation    : X=(A1|A2)&B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA21_4
  CLASS CORE ;
  FOREIGN MDN_OA21_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.18 4.365 0.66 4.595 ;
      RECT  0.43 4.595 0.66 5.46 ;
      RECT  -0.17 5.46 0.66 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.445 1.005 2.06 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.96 1.565 7.955 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  3.96 3.245 7.955 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  3.75 0.6 3.98 1.005 ;
      RECT  3.245 1.005 3.98 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  0.18 1.565 3.475 1.795 ;
      RECT  1.005 1.795 1.235 3.49 ;
      RECT  0.95 0.445 2.705 0.675 ;
      RECT  2.475 0.675 2.705 1.29 ;
      RECT  4.925 2.355 5.155 2.69 ;
      RECT  4.925 2.69 7.395 2.92 ;
      RECT  6.045 2.355 6.275 2.69 ;
      RECT  7.165 2.355 7.395 2.69 ;
      RECT  1.72 4.365 2.76 4.595 ;
  END
END MDN_OA21_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OA21_6
#      Description : One 2-input OR into 2-input AND
#      Equation    : X=(A1|A2)&B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA21_6
  CLASS CORE ;
  FOREIGN MDN_OA21_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 0.98 7.98 1.26 ;
      RECT  7.7 1.26 7.98 1.54 ;
      RECT  7.7 1.54 13.26 1.82 ;
      RECT  11.06 1.82 11.34 3.22 ;
      RECT  7.7 3.22 13.26 3.5 ;
      RECT  7.7 3.5 7.98 4.34 ;
      RECT  6.9 4.34 7.98 4.62 ;
    END
    ANTENNADIFFAREA 9.072 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  10.47 0.37 11.93 0.6 ;
      RECT  4.07 0.445 5.77 0.675 ;
      RECT  4.07 0.675 4.3 1.005 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  4.66 1.005 6.54 1.235 ;
      RECT  6.31 1.235 6.54 1.565 ;
      RECT  6.31 1.565 7.395 1.795 ;
      RECT  7.165 1.795 7.395 2.685 ;
      RECT  7.165 2.685 10.755 2.915 ;
      RECT  8.285 2.355 8.515 2.685 ;
      RECT  9.405 2.355 9.635 2.685 ;
      RECT  10.525 2.355 10.755 2.685 ;
      RECT  7.165 2.915 7.395 3.805 ;
      RECT  6.045 3.805 7.395 4.035 ;
      RECT  6.045 4.035 6.275 4.365 ;
      RECT  2.42 4.365 6.275 4.595 ;
      RECT  11.645 2.35 11.875 2.685 ;
      RECT  11.645 2.685 12.995 2.915 ;
      RECT  12.765 2.35 12.995 2.685 ;
      RECT  0.95 4.925 3.53 5.155 ;
  END
END MDN_OA21_6
#-----------------------------------------------------------------------
#      Cell        : MDN_OA21B_1
#      Description : One 2-input NOR into 2-input NOR
#      Equation    : X=(A1|A2)&!B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA21B_1
  CLASS CORE ;
  FOREIGN MDN_OA21B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 4.65 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 4.3 1.235 ;
      RECT  2.685 1.235 2.915 4.365 ;
      RECT  2.42 4.365 2.915 4.595 ;
    END
    ANTENNADIFFAREA 2.126 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.565 0.37 2.97 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 3.805 ;
      RECT  1.72 3.805 2.355 4.035 ;
  END
END MDN_OA21B_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OA21B_2
#      Description : One 2-input NOR into 2-input NOR
#      Equation    : X=(A1|A2)&!B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA21B_2
  CLASS CORE ;
  FOREIGN MDN_OA21B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.365 1.005 6.54 1.235 ;
      RECT  4.365 1.235 4.595 1.565 ;
      RECT  2.42 1.565 4.595 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  2.42 3.245 4.595 3.475 ;
    END
    ANTENNADIFFAREA 4.252 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.685 ;
      RECT  1.565 2.685 4.035 2.915 ;
      RECT  2.685 2.35 2.915 2.685 ;
      RECT  3.805 2.35 4.035 2.685 ;
      RECT  1.775 2.915 2.005 3.45 ;
      RECT  4.365 4.365 6.54 4.595 ;
      RECT  4.365 4.595 4.595 4.925 ;
      RECT  3.19 4.925 4.595 5.155 ;
  END
END MDN_OA21B_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OA21B_3
#      Description : One 2-input NOR into 2-input NOR
#      Equation    : X=(A1|A2)&!B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA21B_3
  CLASS CORE ;
  FOREIGN MDN_OA21B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 8.54 2.355 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 4.365 8.78 4.595 ;
      RECT  8.285 4.595 8.515 5.46 ;
      RECT  7.84 5.46 9.13 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 8.78 1.235 ;
      RECT  5.485 1.235 5.715 3.245 ;
      RECT  3.19 3.245 5.715 3.475 ;
    END
    ANTENNADIFFAREA 6.054 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 2.685 ;
      RECT  2.685 2.685 5.155 2.915 ;
      RECT  3.805 2.35 4.035 2.685 ;
      RECT  4.925 2.35 5.155 2.685 ;
      RECT  2.685 2.915 2.915 3.805 ;
      RECT  1.72 3.805 2.915 4.035 ;
      RECT  2.42 4.365 4.595 4.595 ;
      RECT  4.365 4.595 4.595 4.925 ;
      RECT  4.365 4.925 8.01 5.155 ;
  END
END MDN_OA21B_3
#-----------------------------------------------------------------------
#      Cell        : MDN_OA21B_4
#      Description : One 2-input NOR into 2-input NOR
#      Equation    : X=(A1|A2)&!B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA21B_4
  CLASS CORE ;
  FOREIGN MDN_OA21B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 10.78 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 11.02 1.235 ;
      RECT  6.605 1.235 6.835 3.245 ;
      RECT  3.19 3.245 6.835 3.475 ;
    END
    ANTENNADIFFAREA 8.18 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 2.685 ;
      RECT  2.685 2.685 6.275 2.915 ;
      RECT  3.805 2.35 4.035 2.685 ;
      RECT  4.925 2.35 5.155 2.685 ;
      RECT  6.045 2.35 6.275 2.685 ;
      RECT  2.685 2.915 2.915 3.805 ;
      RECT  1.72 3.805 2.915 4.035 ;
      RECT  6.605 4.365 11.02 4.595 ;
      RECT  6.605 4.595 6.835 4.925 ;
      RECT  2.42 4.365 4.595 4.595 ;
      RECT  4.365 4.595 4.595 4.925 ;
      RECT  4.365 4.925 6.835 5.155 ;
  END
END MDN_OA21B_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OA221_1
#      Description : Two 2-input ORs into 3-input AND
#      Equation    : X=(A1|A2)&(B1|B2)&C
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA221_1
  CLASS CORE ;
  FOREIGN MDN_OA221_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  1.005 5.46 1.68 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 1.795 0.675 ;
      RECT  1.565 0.675 1.795 1.005 ;
      RECT  1.565 1.005 2.76 1.235 ;
      RECT  1.72 1.565 5.0 1.795 ;
      RECT  1.72 3.805 2.35 4.035 ;
      RECT  2.12 4.035 2.35 4.365 ;
      RECT  2.12 4.365 2.76 4.595 ;
      RECT  4.365 3.805 5.0 4.035 ;
      RECT  4.365 4.035 4.595 4.365 ;
      RECT  3.96 4.365 4.595 4.595 ;
      RECT  4.925 4.365 6.33 4.595 ;
      RECT  4.925 4.595 5.155 4.925 ;
      RECT  6.1 4.595 6.33 5.0 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 1.795 4.595 ;
      RECT  1.565 4.595 1.795 4.925 ;
      RECT  1.565 4.925 5.155 5.155 ;
      RECT  5.99 5.0 6.33 5.23 ;
  END
END MDN_OA221_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OA221_2
#      Description : Two 2-input ORs into 3-input AND
#      Equation    : X=(A1|A2)&(B1|B2)&C
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA221_2
  CLASS CORE ;
  FOREIGN MDN_OA221_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  3.805 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  6.2 3.245 7.24 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 1.795 0.675 ;
      RECT  1.565 0.675 1.795 1.005 ;
      RECT  1.565 1.005 2.76 1.235 ;
      RECT  0.175 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 6.22 4.595 ;
      RECT  5.99 4.595 6.22 5.0 ;
      RECT  5.99 5.0 7.45 5.23 ;
      RECT  1.72 1.565 5.0 1.795 ;
      RECT  1.72 3.805 2.76 4.035 ;
      RECT  3.96 3.805 5.005 4.035 ;
  END
END MDN_OA221_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OA221_4
#      Description : Two 2-input ORs into 3-input AND
#      Equation    : X=(A1|A2)&(B1|B2)&C
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA221_4
  CLASS CORE ;
  FOREIGN MDN_OA221_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.36 -0.14 4.035 0.14 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 9.48 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  6.2 3.245 9.48 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 1.795 0.675 ;
      RECT  1.565 0.675 1.795 1.005 ;
      RECT  1.565 1.005 2.76 1.235 ;
      RECT  1.72 1.565 5.005 1.795 ;
      RECT  8.23 2.41 9.69 2.64 ;
      RECT  1.72 3.805 2.76 4.035 ;
      RECT  3.96 3.805 5.0 4.035 ;
      RECT  7.22 4.365 8.46 4.595 ;
      RECT  7.22 4.595 7.45 5.0 ;
      RECT  8.23 4.595 8.46 5.0 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 6.22 4.595 ;
      RECT  5.99 4.595 6.22 5.0 ;
      RECT  5.99 5.0 7.45 5.23 ;
      RECT  8.23 5.0 8.57 5.23 ;
  END
END MDN_OA221_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OA22_1
#      Description : Two 2-input ORs into 2-input AND
#      Equation    : X=(A1|A2)&(B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA22_1
  CLASS CORE ;
  FOREIGN MDN_OA22_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.96 4.365 5.0 4.595 ;
      RECT  4.365 4.595 4.595 5.46 ;
      RECT  3.92 5.46 5.04 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 5.155 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  4.925 0.14 5.155 1.005 ;
      RECT  4.66 1.005 5.155 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 0.95 5.715 3.53 ;
    END
    ANTENNADIFFAREA 2.566 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 2.65 0.675 ;
      RECT  2.42 0.675 2.65 1.005 ;
      RECT  2.42 1.005 4.3 1.235 ;
      RECT  0.18 1.005 2.06 1.235 ;
      RECT  1.83 1.235 2.06 1.565 ;
      RECT  1.83 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 2.69 ;
      RECT  2.125 1.795 2.355 3.245 ;
      RECT  1.72 3.245 2.76 3.475 ;
  END
END MDN_OA22_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OA22_2
#      Description : Two 2-input ORs into 2-input AND
#      Equation    : X=(A1|A2)&(B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA22_2
  CLASS CORE ;
  FOREIGN MDN_OA22_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 5.715 5.74 ;
      RECT  5.485 4.905 5.715 5.46 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  4.31 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  1.005 -0.14 2.41 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 6.54 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  4.66 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  2.685 1.005 6.22 1.235 ;
      RECT  2.685 1.235 2.915 1.565 ;
      RECT  2.125 1.565 2.915 1.795 ;
      RECT  2.125 1.795 2.355 3.245 ;
      RECT  1.72 3.245 2.76 3.475 ;
      RECT  2.125 0.445 3.53 0.675 ;
      RECT  2.125 0.675 2.355 1.005 ;
      RECT  0.18 1.005 2.355 1.235 ;
  END
END MDN_OA22_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OA22_3
#      Description : Two 2-input ORs into 2-input AND
#      Equation    : X=(A1|A2)&(B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA22_3
  CLASS CORE ;
  FOREIGN MDN_OA22_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 5.715 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  1.005 -0.14 2.41 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 7.24 1.795 ;
      RECT  6.045 1.795 6.275 3.245 ;
      RECT  4.66 3.245 7.24 3.475 ;
    END
    ANTENNADIFFAREA 4.536 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  2.68 1.005 6.22 1.235 ;
      RECT  2.68 1.235 2.91 1.565 ;
      RECT  2.125 1.565 2.91 1.795 ;
      RECT  2.125 1.795 2.355 3.245 ;
      RECT  1.72 3.245 2.76 3.475 ;
      RECT  1.83 0.445 3.53 0.675 ;
      RECT  1.83 0.675 2.06 1.005 ;
      RECT  0.18 1.005 2.06 1.235 ;
  END
END MDN_OA22_3
#-----------------------------------------------------------------------
#      Cell        : MDN_OA22_4
#      Description : Two 2-input ORs into 2-input AND
#      Equation    : X=(A1|A2)&(B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA22_4
  CLASS CORE ;
  FOREIGN MDN_OA22_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 5.715 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  0.0 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  1.005 -0.14 2.41 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 8.78 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  4.66 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 8.57 0.6 ;
      RECT  8.23 0.6 8.46 1.0 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  7.22 0.6 7.45 1.0 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  7.22 1.0 8.46 1.23 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  2.67 1.005 6.22 1.235 ;
      RECT  2.67 1.235 2.9 1.565 ;
      RECT  2.125 1.565 2.9 1.795 ;
      RECT  2.125 1.795 2.355 3.805 ;
      RECT  1.72 3.805 2.76 4.035 ;
      RECT  1.83 0.445 3.53 0.675 ;
      RECT  1.83 0.675 2.06 1.005 ;
      RECT  0.18 1.005 2.06 1.235 ;
  END
END MDN_OA22_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OA22_6
#      Description : Two 2-input ORs into 2-input AND
#      Equation    : X=(A1|A2)&(B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA22_6
  CLASS CORE ;
  FOREIGN MDN_OA22_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.14 0.965 15.5 1.245 ;
      RECT  12.18 1.245 12.46 3.215 ;
      RECT  9.14 3.215 15.5 3.495 ;
    END
    ANTENNADIFFAREA 9.072 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  4.07 0.445 8.01 0.675 ;
      RECT  4.07 0.675 4.3 1.005 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  4.925 1.005 8.515 1.235 ;
      RECT  4.925 1.235 5.155 1.565 ;
      RECT  8.285 1.235 8.515 1.565 ;
      RECT  4.365 1.565 5.155 1.795 ;
      RECT  8.285 1.565 9.635 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  9.405 1.795 9.635 2.685 ;
      RECT  9.405 2.685 11.875 2.915 ;
      RECT  10.525 2.35 10.755 2.685 ;
      RECT  11.645 2.35 11.875 2.685 ;
      RECT  3.19 3.245 5.77 3.475 ;
      RECT  12.765 2.35 12.995 2.685 ;
      RECT  12.765 2.685 15.235 2.915 ;
      RECT  13.885 2.35 14.115 2.685 ;
      RECT  15.005 2.35 15.235 2.685 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.66 4.365 8.78 4.595 ;
      RECT  11.7 4.365 12.94 4.595 ;
      RECT  11.7 4.595 11.93 5.0 ;
      RECT  12.71 4.595 12.94 5.0 ;
      RECT  11.59 5.0 11.93 5.23 ;
      RECT  12.71 5.0 13.05 5.23 ;
  END
END MDN_OA22_6
#-----------------------------------------------------------------------
#      Cell        : MDN_OA2BB2_1
#      Description : One 2-input OR with inverted inputs + 2-input OR into 2-input AND
#      Equation    : X=(!A1|!A2)&(B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA2BB2_1
  CLASS CORE ;
  FOREIGN MDN_OA2BB2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  2.685 4.365 4.3 4.595 ;
      RECT  2.685 4.595 2.915 5.46 ;
      RECT  2.685 5.46 5.715 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  0.0 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      RECT  3.245 0.14 3.475 1.005 ;
      RECT  2.42 1.005 3.475 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.685 1.565 3.53 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  2.42 3.245 2.915 3.475 ;
    END
    ANTENNADIFFAREA 1.992 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.565 0.37 2.97 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  3.96 1.005 5.0 1.235 ;
      RECT  4.66 4.365 5.155 4.595 ;
      RECT  4.925 4.595 5.155 4.925 ;
      RECT  3.19 4.925 5.155 5.155 ;
  END
END MDN_OA2BB2_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OA2BB2_2
#      Description : One 2-input OR with inverted inputs + 2-input OR into 2-input AND
#      Equation    : X=(!A1|!A2)&(B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA2BB2_2
  CLASS CORE ;
  FOREIGN MDN_OA2BB2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 7.42 2.685 ;
      RECT  7.14 2.685 8.54 2.915 ;
      RECT  8.26 2.125 8.54 2.685 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  0.0 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 6.54 1.235 ;
      RECT  4.365 1.235 4.595 3.245 ;
      RECT  2.42 3.245 4.595 3.475 ;
    END
    ANTENNADIFFAREA 4.252 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.445 7.13 0.675 ;
      RECT  6.9 0.675 7.13 1.005 ;
      RECT  6.9 1.005 8.78 1.235 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.685 ;
      RECT  1.565 2.685 4.035 2.915 ;
      RECT  2.685 2.35 2.915 2.685 ;
      RECT  3.805 2.35 4.035 2.685 ;
      RECT  1.565 2.915 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  3.19 4.365 8.78 4.595 ;
  END
END MDN_OA2BB2_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OA2BB2_4
#      Description : One 2-input OR with inverted inputs + 2-input OR into 2-input AND
#      Equation    : X=(!A1|!A2)&(B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA2BB2_4
  CLASS CORE ;
  FOREIGN MDN_OA2BB2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 7.42 2.685 ;
      RECT  7.14 2.685 10.78 2.915 ;
      RECT  8.26 2.125 8.54 2.685 ;
      RECT  9.38 2.125 9.66 2.685 ;
      RECT  10.5 2.125 10.78 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 2.125 15.26 2.355 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 11.02 1.235 ;
      RECT  6.605 1.235 6.835 3.245 ;
      RECT  2.42 3.245 6.835 3.475 ;
    END
    ANTENNADIFFAREA 8.504 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  7.67 0.445 11.61 0.675 ;
      RECT  11.38 0.675 11.61 1.005 ;
      RECT  11.38 1.005 15.5 1.235 ;
      RECT  0.18 1.005 2.06 1.235 ;
      RECT  1.565 1.235 1.795 2.685 ;
      RECT  1.565 2.685 6.275 2.915 ;
      RECT  2.685 2.35 2.915 2.685 ;
      RECT  3.805 2.35 4.035 2.685 ;
      RECT  4.925 2.35 5.155 2.685 ;
      RECT  6.045 2.35 6.275 2.685 ;
      RECT  1.775 2.915 2.005 3.53 ;
      RECT  3.19 4.365 15.5 4.595 ;
  END
END MDN_OA2BB2_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OA311_1
#      Description : One 3-input OR into 3-input AND
#      Equation    : X=(A1|A2|A3)&B1&B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA311_1
  CLASS CORE ;
  FOREIGN MDN_OA311_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  1.005 5.46 1.68 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 6.89 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 6.22 4.595 ;
      RECT  5.99 4.595 6.22 5.0 ;
      RECT  5.99 5.0 6.33 5.23 ;
      RECT  1.72 1.005 5.0 1.235 ;
      RECT  3.96 3.805 5.0 4.035 ;
  END
END MDN_OA311_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OA311_2
#      Description : One 3-input OR into 3-input AND
#      Equation    : X=(A1|A2|A3)&B1&B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA311_2
  CLASS CORE ;
  FOREIGN MDN_OA311_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 0.14 3.475 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  6.2 3.245 7.24 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 6.22 4.595 ;
      RECT  5.99 4.595 6.22 5.0 ;
      RECT  5.99 5.0 7.45 5.23 ;
      RECT  1.72 1.005 5.0 1.235 ;
      RECT  3.96 3.805 5.0 4.035 ;
  END
END MDN_OA311_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OA311_4
#      Description : One 3-input OR into 3-input AND
#      Equation    : X=(A1|A2|A3)&B1&B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA311_4
  CLASS CORE ;
  FOREIGN MDN_OA311_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 9.48 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  6.2 3.245 9.48 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.005 5.0 1.235 ;
      RECT  8.23 2.4 9.69 2.63 ;
      RECT  3.96 3.805 5.0 4.035 ;
      RECT  7.22 4.365 8.46 4.595 ;
      RECT  7.22 4.595 7.45 5.0 ;
      RECT  8.23 4.595 8.46 5.0 ;
      RECT  0.18 1.005 1.235 1.235 ;
      RECT  1.005 1.235 1.235 4.365 ;
      RECT  0.18 4.365 6.22 4.595 ;
      RECT  5.99 4.595 6.22 5.0 ;
      RECT  5.99 5.0 7.45 5.23 ;
      RECT  8.23 5.0 8.57 5.23 ;
  END
END MDN_OA311_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OA31_1
#      Description : One 3-input OR into 2-input AND
#      Equation    : X=(A1|A2|A3)&B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA31_1
  CLASS CORE ;
  FOREIGN MDN_OA31_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.89 5.74 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 4.48 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  0.0 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.36 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.705 0.14 3.935 1.005 ;
      RECT  2.42 1.005 3.935 1.235 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 3.245 ;
      RECT  4.66 3.245 5.155 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  4.195 0.37 5.21 0.6 ;
      RECT  4.195 0.6 4.425 1.565 ;
      RECT  3.245 1.565 4.425 1.795 ;
      RECT  3.245 1.795 3.475 3.5 ;
      RECT  1.835 0.435 3.475 0.665 ;
      RECT  3.245 0.665 3.475 0.775 ;
      RECT  1.835 0.665 2.065 1.005 ;
      RECT  0.18 1.005 2.065 1.235 ;
      RECT  1.72 4.365 2.76 4.595 ;
  END
END MDN_OA31_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OA31_2
#      Description : One 3-input OR into 2-input AND
#      Equation    : X=(A1|A2|A3)&B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA31_2
  CLASS CORE ;
  FOREIGN MDN_OA31_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 5.715 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  0.0 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.36 -0.14 3.99 0.14 ;
      RECT  3.76 0.14 3.99 1.005 ;
      RECT  2.42 1.005 3.99 1.235 ;
      RECT  1.005 -0.14 2.41 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 6.54 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  4.66 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  4.555 1.005 6.22 1.01 ;
      RECT  4.55 1.01 6.22 1.015 ;
      RECT  4.545 1.015 6.22 1.02 ;
      RECT  4.54 1.02 6.22 1.025 ;
      RECT  4.535 1.025 6.22 1.03 ;
      RECT  4.53 1.03 6.22 1.035 ;
      RECT  4.525 1.035 6.22 1.04 ;
      RECT  4.52 1.04 6.22 1.045 ;
      RECT  4.515 1.045 6.22 1.05 ;
      RECT  4.51 1.05 6.22 1.055 ;
      RECT  4.505 1.055 6.22 1.06 ;
      RECT  4.5 1.06 6.22 1.065 ;
      RECT  4.495 1.065 6.22 1.07 ;
      RECT  4.49 1.07 6.22 1.075 ;
      RECT  4.485 1.075 6.22 1.08 ;
      RECT  4.48 1.08 6.22 1.085 ;
      RECT  4.475 1.085 6.22 1.09 ;
      RECT  4.47 1.09 6.22 1.095 ;
      RECT  4.465 1.095 6.22 1.1 ;
      RECT  4.46 1.1 6.22 1.105 ;
      RECT  4.455 1.105 6.22 1.11 ;
      RECT  4.45 1.11 6.22 1.115 ;
      RECT  4.445 1.115 6.22 1.12 ;
      RECT  4.44 1.12 6.22 1.125 ;
      RECT  4.435 1.125 6.22 1.13 ;
      RECT  4.43 1.13 6.22 1.135 ;
      RECT  4.425 1.135 6.22 1.14 ;
      RECT  4.42 1.14 6.22 1.145 ;
      RECT  4.415 1.145 6.22 1.15 ;
      RECT  4.41 1.15 6.22 1.155 ;
      RECT  4.405 1.155 6.22 1.16 ;
      RECT  4.4 1.16 6.22 1.165 ;
      RECT  4.395 1.165 6.22 1.17 ;
      RECT  4.39 1.17 6.22 1.175 ;
      RECT  4.385 1.175 6.22 1.18 ;
      RECT  4.38 1.18 6.22 1.185 ;
      RECT  4.375 1.185 6.22 1.19 ;
      RECT  4.37 1.19 6.22 1.195 ;
      RECT  4.365 1.195 6.22 1.2 ;
      RECT  4.36 1.2 6.22 1.205 ;
      RECT  4.355 1.205 6.22 1.21 ;
      RECT  4.35 1.21 6.22 1.215 ;
      RECT  4.345 1.215 6.22 1.22 ;
      RECT  4.34 1.22 6.22 1.225 ;
      RECT  4.335 1.225 6.22 1.23 ;
      RECT  4.33 1.23 6.22 1.235 ;
      RECT  4.325 1.235 4.65 1.24 ;
      RECT  4.32 1.24 4.645 1.245 ;
      RECT  4.315 1.245 4.64 1.25 ;
      RECT  4.31 1.25 4.635 1.255 ;
      RECT  4.305 1.255 4.63 1.26 ;
      RECT  4.3 1.26 4.625 1.265 ;
      RECT  4.295 1.265 4.62 1.27 ;
      RECT  4.29 1.27 4.615 1.275 ;
      RECT  4.285 1.275 4.61 1.28 ;
      RECT  4.28 1.28 4.605 1.285 ;
      RECT  4.275 1.285 4.6 1.29 ;
      RECT  4.27 1.29 4.595 1.295 ;
      RECT  4.265 1.295 4.59 1.3 ;
      RECT  4.26 1.3 4.585 1.305 ;
      RECT  4.255 1.305 4.58 1.31 ;
      RECT  4.25 1.31 4.575 1.315 ;
      RECT  4.245 1.315 4.57 1.32 ;
      RECT  4.24 1.32 4.565 1.325 ;
      RECT  4.235 1.325 4.56 1.33 ;
      RECT  4.23 1.33 4.555 1.335 ;
      RECT  4.225 1.335 4.55 1.34 ;
      RECT  4.22 1.34 4.545 1.345 ;
      RECT  4.215 1.345 4.54 1.35 ;
      RECT  4.21 1.35 4.535 1.355 ;
      RECT  4.205 1.355 4.53 1.36 ;
      RECT  4.2 1.36 4.525 1.365 ;
      RECT  4.195 1.365 4.52 1.37 ;
      RECT  4.19 1.37 4.515 1.375 ;
      RECT  4.185 1.375 4.51 1.38 ;
      RECT  4.18 1.38 4.505 1.385 ;
      RECT  4.175 1.385 4.5 1.39 ;
      RECT  4.17 1.39 4.495 1.395 ;
      RECT  4.165 1.395 4.49 1.4 ;
      RECT  4.16 1.4 4.485 1.405 ;
      RECT  4.155 1.405 4.48 1.41 ;
      RECT  4.15 1.41 4.475 1.415 ;
      RECT  4.145 1.415 4.47 1.42 ;
      RECT  4.14 1.42 4.465 1.425 ;
      RECT  4.135 1.425 4.46 1.43 ;
      RECT  4.13 1.43 4.455 1.435 ;
      RECT  4.125 1.435 4.45 1.44 ;
      RECT  4.12 1.44 4.445 1.445 ;
      RECT  4.115 1.445 4.44 1.45 ;
      RECT  4.11 1.45 4.435 1.455 ;
      RECT  4.105 1.455 4.43 1.46 ;
      RECT  4.1 1.46 4.425 1.465 ;
      RECT  4.095 1.465 4.42 1.47 ;
      RECT  4.09 1.47 4.415 1.475 ;
      RECT  4.085 1.475 4.41 1.48 ;
      RECT  4.08 1.48 4.405 1.485 ;
      RECT  4.075 1.485 4.4 1.49 ;
      RECT  4.07 1.49 4.395 1.495 ;
      RECT  4.07 1.495 4.39 1.5 ;
      RECT  4.07 1.5 4.385 1.505 ;
      RECT  4.07 1.505 4.38 1.51 ;
      RECT  4.07 1.51 4.375 1.515 ;
      RECT  4.07 1.515 4.37 1.52 ;
      RECT  4.07 1.52 4.365 1.525 ;
      RECT  4.07 1.525 4.36 1.53 ;
      RECT  4.07 1.53 4.355 1.535 ;
      RECT  4.07 1.535 4.35 1.54 ;
      RECT  4.07 1.54 4.345 1.545 ;
      RECT  4.07 1.545 4.34 1.55 ;
      RECT  4.07 1.55 4.335 1.555 ;
      RECT  4.07 1.555 4.33 1.56 ;
      RECT  4.07 1.56 4.325 1.565 ;
      RECT  3.245 1.565 4.32 1.57 ;
      RECT  3.245 1.57 4.315 1.575 ;
      RECT  3.245 1.575 4.31 1.58 ;
      RECT  3.245 1.58 4.305 1.585 ;
      RECT  3.245 1.585 4.3 1.795 ;
      RECT  3.245 1.795 3.475 3.53 ;
      RECT  1.83 0.445 3.53 0.675 ;
      RECT  1.83 0.675 2.06 1.005 ;
      RECT  0.18 1.005 2.06 1.235 ;
      RECT  1.72 4.365 2.765 4.595 ;
  END
END MDN_OA31_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OA31_4
#      Description : One 3-input OR into 2-input AND
#      Equation    : X=(A1|A2|A3)&B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA31_4
  CLASS CORE ;
  FOREIGN MDN_OA31_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 5.715 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  0.0 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.36 -0.14 3.99 0.14 ;
      RECT  3.76 0.14 3.99 1.005 ;
      RECT  2.42 1.005 3.99 1.235 ;
      RECT  1.005 -0.14 2.41 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.715 1.565 8.78 1.795 ;
      RECT  4.715 1.795 4.945 1.905 ;
      RECT  6.6 1.795 6.83 3.245 ;
      RECT  4.66 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  4.255 1.005 6.22 1.235 ;
      RECT  4.255 1.235 4.485 1.565 ;
      RECT  3.245 1.565 4.485 1.795 ;
      RECT  3.245 1.795 3.475 3.5 ;
      RECT  1.83 0.445 3.53 0.675 ;
      RECT  1.83 0.675 2.06 1.005 ;
      RECT  0.18 1.005 2.06 1.235 ;
      RECT  7.325 2.35 7.555 2.685 ;
      RECT  7.32 2.685 8.515 2.915 ;
      RECT  8.285 2.35 8.515 2.685 ;
      RECT  1.72 4.365 2.76 4.595 ;
  END
END MDN_OA31_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OA32_1
#      Description : One 3-input OR + one 2-input OR into 2-input AND
#      Equation    : X=(A1|A2|A3)&(B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA32_1
  CLASS CORE ;
  FOREIGN MDN_OA32_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  5.485 0.14 5.715 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  5.485 1.005 6.22 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 5.715 1.795 ;
      RECT  2.125 1.795 2.355 3.805 ;
      RECT  1.72 3.805 2.76 4.035 ;
      RECT  0.95 0.445 2.355 0.675 ;
      RECT  2.125 0.675 2.355 1.005 ;
      RECT  2.125 1.005 5.0 1.235 ;
      RECT  3.96 4.365 5.0 4.595 ;
  END
END MDN_OA32_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OA32_2
#      Description : One 3-input OR + one 2-input OR into 2-input AND
#      Equation    : X=(A1|A2|A3)&(B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA32_2
  CLASS CORE ;
  FOREIGN MDN_OA32_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  4.31 5.46 5.715 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  0.0 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  5.485 0.14 5.715 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  6.2 3.245 7.24 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  5.485 1.005 6.22 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 5.715 1.795 ;
      RECT  2.125 1.795 2.355 3.805 ;
      RECT  1.72 3.805 2.76 4.035 ;
      RECT  0.95 0.445 2.355 0.675 ;
      RECT  2.125 0.675 2.355 1.005 ;
      RECT  2.125 1.005 5.0 1.235 ;
      RECT  3.96 4.365 5.0 4.595 ;
  END
END MDN_OA32_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OA32_4
#      Description : One 3-input OR + one 2-input OR into 2-input AND
#      Equation    : X=(A1|A2|A3)&(B1|B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA32_4
  CLASS CORE ;
  FOREIGN MDN_OA32_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 9.48 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  6.2 3.245 9.48 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 9.69 0.6 ;
      RECT  8.23 0.6 8.46 1.005 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  7.22 0.6 7.45 1.005 ;
      RECT  5.485 1.005 6.22 1.235 ;
      RECT  7.22 1.005 8.46 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 5.715 1.795 ;
      RECT  2.125 1.795 2.355 3.805 ;
      RECT  1.72 3.805 2.76 4.035 ;
      RECT  0.95 0.445 2.355 0.675 ;
      RECT  2.125 0.675 2.355 1.005 ;
      RECT  2.125 1.005 5.0 1.235 ;
      RECT  3.96 4.365 5.0 4.595 ;
  END
END MDN_OA32_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OA41_1
#      Description : One 4-input OR into 2-input AND
#      Equation    : X=(A1|A2|A3|A4)&B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA41_1
  CLASS CORE ;
  FOREIGN MDN_OA41_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A4
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.445 1.005 2.06 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 1.565 6.54 1.795 ;
      RECT  6.045 1.795 6.275 3.245 ;
      RECT  6.045 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  5.485 1.005 6.22 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  0.18 1.565 5.715 1.795 ;
      RECT  1.005 1.795 1.235 3.5 ;
      RECT  0.95 0.445 2.65 0.675 ;
      RECT  2.42 0.675 2.65 1.005 ;
      RECT  2.42 1.005 5.0 1.235 ;
      RECT  1.72 4.365 2.76 4.595 ;
      RECT  3.96 4.365 5.0 4.595 ;
  END
END MDN_OA41_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OA41_2
#      Description : One 4-input OR into 2-input AND
#      Equation    : X=(A1|A2|A3|A4)&B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA41_2
  CLASS CORE ;
  FOREIGN MDN_OA41_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 4.365 2.94 5.0 ;
      RECT  2.63 5.0 2.97 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A4
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.35 0.7 3.475 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 9.13 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  1.565 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  1.565 0.14 1.795 0.935 ;
      RECT  1.565 0.935 2.06 1.165 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 7.24 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  6.2 3.245 7.24 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  5.485 1.005 6.22 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  3.245 1.565 5.715 1.795 ;
      RECT  3.245 1.795 3.475 2.125 ;
      RECT  0.18 1.565 0.675 1.795 ;
      RECT  0.445 1.795 0.675 1.855 ;
      RECT  0.445 1.855 1.235 2.085 ;
      RECT  1.005 2.085 1.235 2.125 ;
      RECT  1.005 2.125 3.475 2.355 ;
      RECT  3.245 2.355 3.475 2.36 ;
      RECT  1.005 2.355 1.235 3.53 ;
      RECT  2.42 1.005 5.0 1.235 ;
      RECT  2.42 1.235 2.65 1.395 ;
      RECT  0.95 1.395 2.65 1.625 ;
      RECT  1.72 3.245 2.76 3.475 ;
      RECT  3.96 4.365 5.0 4.595 ;
  END
END MDN_OA41_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OA41_4
#      Description : One 4-input OR into 2-input AND
#      Equation    : X=(A1|A2|A3|A4)&B
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OA41_4
  CLASS CORE ;
  FOREIGN MDN_OA41_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 4.365 2.94 5.0 ;
      RECT  2.63 5.0 2.97 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A4
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.35 0.7 3.475 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  1.565 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  1.565 0.14 1.795 0.945 ;
      RECT  1.565 0.945 2.06 1.175 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.2 1.565 9.48 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  6.2 3.245 9.48 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 9.69 0.6 ;
      RECT  8.23 0.6 8.46 1.005 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  7.22 0.6 7.45 1.005 ;
      RECT  5.485 1.005 6.22 1.235 ;
      RECT  7.22 1.005 8.46 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  3.245 1.565 5.715 1.795 ;
      RECT  3.245 1.795 3.475 2.125 ;
      RECT  0.18 1.565 0.675 1.795 ;
      RECT  0.445 1.795 0.675 1.875 ;
      RECT  0.445 1.875 1.235 2.105 ;
      RECT  1.005 2.105 1.235 2.125 ;
      RECT  1.005 2.125 3.475 2.355 ;
      RECT  1.005 2.355 1.235 3.53 ;
      RECT  2.42 1.005 5.0 1.235 ;
      RECT  2.42 1.235 2.65 1.41 ;
      RECT  0.95 1.41 2.65 1.64 ;
      RECT  1.72 3.245 2.76 3.475 ;
      RECT  3.96 4.365 5.0 4.595 ;
  END
END MDN_OA41_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI2111_1
#      Description : One 2-input OR into 4-input NAND
#      Equation    : X=!((A1|A2)&B1&B2&B3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI2111_1
  CLASS CORE ;
  FOREIGN MDN_OAI2111_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 4.48 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  1.005 5.46 2.41 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 -0.14 2.915 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      RECT  2.685 0.14 2.915 1.005 ;
      RECT  2.42 1.005 2.915 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 1.005 6.54 1.235 ;
      RECT  5.485 1.235 5.715 1.565 ;
      RECT  4.365 1.565 5.715 1.795 ;
      RECT  4.365 1.795 4.595 3.805 ;
      RECT  3.19 3.805 5.155 4.035 ;
      RECT  4.925 4.035 5.155 4.365 ;
      RECT  4.925 4.365 6.54 4.595 ;
    END
    ANTENNADIFFAREA 3.882 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.96 1.005 5.0 1.235 ;
      RECT  1.72 1.565 3.53 1.795 ;
      RECT  1.72 4.365 2.76 4.595 ;
  END
END MDN_OAI2111_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI2111_2
#      Description : One 2-input OR into 4-input NAND
#      Equation    : X=!((A1|A2)&B1&B2&B3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI2111_2
  CLASS CORE ;
  FOREIGN MDN_OAI2111_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 10.78 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 -0.14 11.37 0.14 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.405 1.005 11.02 1.235 ;
      RECT  9.405 1.235 9.635 1.565 ;
      RECT  8.845 1.565 9.635 1.795 ;
      RECT  8.845 1.795 9.075 4.365 ;
      RECT  2.42 4.365 11.02 4.595 ;
    END
    ANTENNADIFFAREA 8.412 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.445 7.13 0.675 ;
      RECT  6.9 0.675 7.13 1.005 ;
      RECT  6.9 1.005 8.78 1.235 ;
      RECT  7.67 0.445 10.25 0.675 ;
      RECT  0.18 1.005 6.54 1.235 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  1.83 4.595 2.06 4.925 ;
      RECT  1.83 4.925 3.53 5.155 ;
  END
END MDN_OAI2111_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI2111_4
#      Description : One 2-input OR into 4-input NAND
#      Equation    : X=!((A1|A2)&B1&B2&B3)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI2111_4
  CLASS CORE ;
  FOREIGN MDN_OAI2111_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.34 2.125 21.98 2.355 ;
      RECT  18.34 2.355 18.62 2.915 ;
      RECT  19.46 2.355 19.74 2.915 ;
      RECT  20.58 2.355 20.86 2.915 ;
      RECT  21.7 2.355 21.98 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.84 -0.14 22.57 0.14 ;
      RECT  10.64 -0.14 11.76 0.14 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.365 1.005 22.22 1.235 ;
      RECT  18.365 1.235 18.595 1.565 ;
      RECT  17.805 1.565 18.595 1.795 ;
      RECT  17.805 1.795 18.035 4.365 ;
      RECT  4.66 4.365 22.22 4.595 ;
    END
    ANTENNADIFFAREA 16.824 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.55 0.445 12.49 0.675 ;
      RECT  8.55 0.675 8.78 1.005 ;
      RECT  0.18 1.005 8.78 1.235 ;
      RECT  14.39 0.445 21.45 0.675 ;
      RECT  9.14 1.005 17.74 1.235 ;
      RECT  0.18 4.365 4.305 4.595 ;
      RECT  4.075 4.595 4.305 4.925 ;
      RECT  4.075 4.925 8.01 5.155 ;
  END
END MDN_OAI2111_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI211_1
#      Description : One 2-input OR into 3-input NAND
#      Equation    : X=!((A1|A2)&B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI211_1
  CLASS CORE ;
  FOREIGN MDN_OAI211_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 1.005 4.3 1.235 ;
      RECT  3.245 1.235 3.475 3.805 ;
      RECT  1.72 3.805 4.3 4.035 ;
    END
    ANTENNADIFFAREA 3.308 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 2.76 1.235 ;
  END
END MDN_OAI211_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI211_2
#      Description : One 2-input OR into 3-input NAND
#      Equation    : X=!((A1|A2)&B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI211_2
  CLASS CORE ;
  FOREIGN MDN_OAI211_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 7.955 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      RECT  3.245 0.14 3.475 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.165 1.005 8.78 1.235 ;
      RECT  7.165 1.235 7.395 1.565 ;
      RECT  6.605 1.565 7.395 1.795 ;
      RECT  6.605 1.795 6.835 4.365 ;
      RECT  2.42 4.365 8.78 4.595 ;
    END
    ANTENNADIFFAREA 6.616 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.445 8.01 0.675 ;
      RECT  0.18 1.005 6.54 1.235 ;
      RECT  0.95 4.925 3.53 5.155 ;
  END
END MDN_OAI211_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI211_3
#      Description : One 2-input OR into 3-input NAND
#      Equation    : X=!((A1|A2)&B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI211_3
  CLASS CORE ;
  FOREIGN MDN_OAI211_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 7.42 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 16.38 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 11.9 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.895 12.435 5.46 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.8 -0.14 18.09 0.14 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.325 1.565 16.97 1.795 ;
      RECT  13.325 1.795 13.555 4.365 ;
      RECT  4.66 4.365 16.2 4.595 ;
    END
    ANTENNADIFFAREA 10.404 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.285 0.445 12.49 0.675 ;
      RECT  8.285 0.675 8.515 1.005 ;
      RECT  0.18 1.005 8.515 1.235 ;
      RECT  12.765 0.445 15.795 0.675 ;
      RECT  12.765 0.675 12.995 1.005 ;
      RECT  15.565 0.675 15.795 1.005 ;
      RECT  9.14 1.005 12.995 1.235 ;
      RECT  15.565 1.005 16.2 1.235 ;
      RECT  0.18 4.365 4.035 4.595 ;
      RECT  3.805 4.595 4.035 4.925 ;
      RECT  3.805 4.925 8.01 5.155 ;
  END
END MDN_OAI211_3
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI211_4
#      Description : One 2-input OR into 3-input NAND
#      Equation    : X=!((A1|A2)&B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI211_4
  CLASS CORE ;
  FOREIGN MDN_OAI211_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.8 -0.14 18.09 0.14 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.325 1.565 17.74 1.795 ;
      RECT  13.325 1.795 13.555 4.365 ;
      RECT  9.14 4.365 17.74 4.595 ;
      RECT  9.14 4.595 9.37 4.925 ;
      RECT  5.43 4.925 9.37 5.155 ;
    END
    ANTENNADIFFAREA 12.584 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.55 0.445 12.49 0.675 ;
      RECT  8.55 0.675 8.78 1.005 ;
      RECT  0.18 1.005 8.78 1.235 ;
      RECT  13.325 0.445 16.97 0.675 ;
      RECT  13.325 0.675 13.555 1.005 ;
      RECT  9.14 1.005 13.555 1.235 ;
      RECT  0.18 4.365 8.78 4.595 ;
  END
END MDN_OAI211_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI21_1
#      Description : One 2-input OR into 2-input NAND
#      Equation    : X=!((A1|A2)&B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI21_1
  CLASS CORE ;
  FOREIGN MDN_OAI21_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.125 1.565 3.53 1.795 ;
      RECT  2.125 1.795 2.355 3.805 ;
      RECT  1.72 3.805 2.76 4.035 ;
    END
    ANTENNADIFFAREA 2.89 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 2.76 1.235 ;
  END
END MDN_OAI21_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI21_2
#      Description : One 2-input OR into 2-input NAND
#      Equation    : X=!((A1|A2)&B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI21_2
  CLASS CORE ;
  FOREIGN MDN_OAI21_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  1.005 5.46 2.41 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      RECT  3.245 0.14 3.475 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.925 1.005 6.54 1.235 ;
      RECT  4.925 1.235 5.155 1.565 ;
      RECT  4.365 1.565 5.155 1.795 ;
      RECT  4.365 1.795 4.595 4.365 ;
      RECT  2.42 4.365 6.54 4.595 ;
    END
    ANTENNADIFFAREA 4.82 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  4.365 0.445 5.77 0.675 ;
      RECT  4.365 0.675 4.595 1.005 ;
      RECT  0.18 1.005 4.595 1.235 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  1.83 4.595 2.06 4.925 ;
      RECT  1.83 4.925 3.53 5.155 ;
  END
END MDN_OAI21_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI21_3
#      Description : One 2-input OR into 2-input NAND
#      Equation    : X=!((A1|A2)&B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI21_3
  CLASS CORE ;
  FOREIGN MDN_OAI21_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 6.3 2.355 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 9.66 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 -0.14 11.37 0.14 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.165 1.005 9.48 1.235 ;
      RECT  7.165 1.235 7.395 1.565 ;
      RECT  6.605 1.565 7.395 1.795 ;
      RECT  6.605 1.795 6.835 3.805 ;
      RECT  3.96 3.805 9.48 4.035 ;
    END
    ANTENNADIFFAREA 7.23 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  6.605 0.445 10.25 0.675 ;
      RECT  6.605 0.675 6.835 1.005 ;
      RECT  0.18 1.005 6.835 1.235 ;
      RECT  0.95 4.925 5.77 5.155 ;
  END
END MDN_OAI21_3
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI21_4
#      Description : One 2-input OR into 2-input NAND
#      Equation    : X=!((A1|A2)&B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI21_4
  CLASS CORE ;
  FOREIGN MDN_OAI21_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.88 -0.14 13.61 0.14 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.405 1.005 13.26 1.235 ;
      RECT  9.405 1.235 9.635 1.565 ;
      RECT  8.845 1.565 9.635 1.795 ;
      RECT  8.845 1.795 9.075 4.365 ;
      RECT  4.66 4.365 13.26 4.595 ;
    END
    ANTENNADIFFAREA 9.64 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.845 0.445 12.49 0.675 ;
      RECT  8.845 0.675 9.075 1.005 ;
      RECT  0.18 1.005 9.075 1.235 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.07 4.595 4.3 4.925 ;
      RECT  4.07 4.925 8.01 5.155 ;
  END
END MDN_OAI21_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI21B_1
#      Description : One 2-input OR into 2-input NAND (other input inverted)
#      Equation    : X=!((A1|A2)&!B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI21B_1
  CLASS CORE ;
  FOREIGN MDN_OAI21B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.365 2.06 4.595 ;
      RECT  1.005 4.595 1.235 5.46 ;
      RECT  1.005 5.46 3.475 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.68 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 1.005 2.06 1.235 ;
      RECT  1.005 1.235 1.235 3.53 ;
    END
    ANTENNADIFFAREA 2.086 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 2.61 0.675 ;
      RECT  2.38 0.675 2.61 1.005 ;
      RECT  2.38 1.005 2.76 1.235 ;
      RECT  3.245 1.005 4.3 1.235 ;
      RECT  3.245 1.235 3.475 4.365 ;
      RECT  2.395 4.365 4.3 4.595 ;
      RECT  2.395 4.595 2.625 4.925 ;
      RECT  1.51 4.925 2.625 5.155 ;
      RECT  1.51 5.155 1.85 5.23 ;
      RECT  0.18 3.805 2.76 4.035 ;
  END
END MDN_OAI21B_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI21B_2
#      Description : One 2-input OR into 2-input NAND (other input inverted)
#      Equation    : X=!((A1|A2)&!B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI21B_2
  CLASS CORE ;
  FOREIGN MDN_OAI21B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.685 ;
      RECT  2.66 2.685 4.06 2.915 ;
      RECT  3.78 2.125 4.06 2.685 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 1.82 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 4.365 7.42 5.0 ;
      RECT  7.11 5.0 7.45 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      RECT  3.245 0.14 3.475 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.365 1.565 6.54 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  2.42 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 4.82 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  4.365 0.445 5.77 0.675 ;
      RECT  4.365 0.675 4.595 1.005 ;
      RECT  0.18 1.005 4.595 1.235 ;
      RECT  6.9 1.565 7.395 1.795 ;
      RECT  7.165 1.795 7.395 2.405 ;
      RECT  4.98 2.405 7.395 2.635 ;
      RECT  7.165 2.635 7.395 3.245 ;
      RECT  6.9 3.245 7.395 3.475 ;
      RECT  0.18 4.365 2.355 4.595 ;
      RECT  2.125 4.595 2.355 4.925 ;
      RECT  2.125 4.925 3.53 5.155 ;
  END
END MDN_OAI21B_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI21B_3
#      Description : One 2-input OR into 2-input NAND (other input inverted)
#      Equation    : X=!((A1|A2)&!B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI21B_3
  CLASS CORE ;
  FOREIGN MDN_OAI21B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.685 ;
      RECT  3.78 2.685 6.3 2.915 ;
      RECT  4.9 2.125 5.18 2.685 ;
      RECT  6.02 2.125 6.3 2.685 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 2.94 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
      RECT  2.66 2.125 2.94 2.685 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 2.125 11.9 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 2.8 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  5.485 -0.14 6.89 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      RECT  3.245 0.14 3.475 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.605 1.565 9.48 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  6.605 3.245 9.48 3.475 ;
      RECT  6.605 3.475 6.835 3.805 ;
      RECT  3.96 3.805 6.835 4.035 ;
    END
    ANTENNADIFFAREA 7.23 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  6.31 0.445 10.25 0.675 ;
      RECT  6.31 0.675 6.54 1.005 ;
      RECT  0.18 1.005 6.54 1.235 ;
      RECT  9.965 1.565 11.72 1.795 ;
      RECT  9.965 1.795 10.195 2.685 ;
      RECT  7.165 2.35 7.395 2.685 ;
      RECT  7.165 2.685 10.195 2.915 ;
      RECT  8.285 2.35 8.515 2.685 ;
      RECT  9.405 2.35 9.635 2.685 ;
      RECT  9.965 2.915 10.195 3.245 ;
      RECT  9.965 3.245 11.72 3.475 ;
      RECT  0.95 4.925 5.77 5.155 ;
  END
END MDN_OAI21B_3
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI21B_4
#      Description : One 2-input OR into 2-input NAND (other input inverted)
#      Equation    : X=!((A1|A2)&!B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI21B_4
  CLASS CORE ;
  FOREIGN MDN_OAI21B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.68 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.685 ;
      RECT  4.9 2.685 8.54 2.915 ;
      RECT  6.02 2.125 6.3 2.685 ;
      RECT  7.14 2.125 7.42 2.685 ;
      RECT  8.26 2.125 8.54 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.685 ;
      RECT  0.42 2.685 4.06 2.915 ;
      RECT  1.54 2.125 1.82 2.685 ;
      RECT  2.66 2.125 2.94 2.685 ;
      RECT  3.78 2.125 4.06 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 4.365 14.14 5.0 ;
      RECT  13.83 5.0 14.17 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.85 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 3.475 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 15.68 5.74 ;
      LAYER VIA12 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 -0.14 15.85 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 15.68 0.14 ;
      LAYER VIA12 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.405 1.005 13.26 1.235 ;
      RECT  9.405 1.235 9.635 1.565 ;
      RECT  8.845 1.565 9.635 1.795 ;
      RECT  8.845 1.795 9.075 3.805 ;
      RECT  4.66 3.805 13.26 4.035 ;
    END
    ANTENNADIFFAREA 9.64 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.845 0.445 12.49 0.675 ;
      RECT  8.845 0.675 9.075 1.005 ;
      RECT  0.18 1.005 9.075 1.235 ;
      RECT  13.62 1.565 14.115 1.795 ;
      RECT  13.885 1.795 14.115 2.685 ;
      RECT  9.38 2.125 9.66 2.685 ;
      RECT  9.38 2.685 14.115 2.915 ;
      RECT  10.5 2.125 10.78 2.685 ;
      RECT  11.62 2.125 11.9 2.685 ;
      RECT  12.74 2.125 13.02 2.685 ;
      RECT  13.885 2.915 14.115 3.245 ;
      RECT  13.62 3.245 14.115 3.475 ;
      RECT  0.18 4.365 8.01 4.595 ;
  END
END MDN_OAI21B_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI221_1
#      Description : Two 2-input ORs into 3-input NAND
#      Equation    : X=!((A1|A2)&(B1|B2)&C)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI221_1
  CLASS CORE ;
  FOREIGN MDN_OAI221_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  1.005 5.46 2.41 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 -0.14 2.915 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      RECT  2.685 0.14 2.915 1.005 ;
      RECT  2.42 1.005 2.915 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.365 1.565 5.0 1.795 ;
      RECT  4.365 1.795 4.595 3.805 ;
      RECT  3.19 3.805 5.0 4.035 ;
    END
    ANTENNADIFFAREA 2.984 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.245 0.445 6.275 0.675 ;
      RECT  6.045 0.675 6.275 1.005 ;
      RECT  3.245 0.675 3.475 1.565 ;
      RECT  6.045 1.005 6.54 1.235 ;
      RECT  1.72 1.565 3.475 1.795 ;
      RECT  3.96 1.005 5.77 1.235 ;
      RECT  1.72 4.365 2.76 4.595 ;
      RECT  3.96 4.365 6.54 4.595 ;
  END
END MDN_OAI221_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI221_2
#      Description : Two 2-input ORs into 3-input NAND
#      Equation    : X=!((A1|A2)&(B1|B2)&C)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI221_2
  CLASS CORE ;
  FOREIGN MDN_OAI221_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 10.78 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.08 -0.14 11.37 0.14 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  5.43 1.565 6.835 1.795 ;
      RECT  6.605 1.795 6.835 4.365 ;
      RECT  2.42 4.365 8.78 4.595 ;
    END
    ANTENNADIFFAREA 6.482 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  4.07 0.445 10.25 0.675 ;
      RECT  4.07 0.675 4.3 1.005 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  4.66 1.005 11.02 1.235 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  1.83 4.595 2.06 4.925 ;
      RECT  1.83 4.925 3.53 5.155 ;
      RECT  9.14 4.365 11.02 4.595 ;
      RECT  9.14 4.595 9.37 4.925 ;
      RECT  7.67 4.925 9.37 5.155 ;
  END
END MDN_OAI221_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI221_4
#      Description : Two 2-input ORs into 3-input NAND
#      Equation    : X=!((A1|A2)&(B1|B2)&C)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI221_4
  CLASS CORE ;
  FOREIGN MDN_OAI221_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.685 ;
      RECT  4.9 2.685 8.54 2.915 ;
      RECT  6.02 2.125 6.3 2.685 ;
      RECT  7.14 2.125 7.42 2.685 ;
      RECT  8.26 2.125 8.54 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 14.14 2.685 ;
      RECT  13.86 2.685 17.5 2.915 ;
      RECT  14.98 2.125 15.26 2.685 ;
      RECT  16.1 2.125 16.38 2.685 ;
      RECT  17.22 2.125 17.5 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.34 2.125 21.98 2.355 ;
      RECT  18.34 2.355 18.62 2.915 ;
      RECT  19.46 2.355 19.74 2.915 ;
      RECT  20.58 2.355 20.86 2.915 ;
      RECT  21.7 2.355 21.98 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.685 ;
      RECT  9.38 2.685 13.02 2.915 ;
      RECT  10.5 2.125 10.78 2.685 ;
      RECT  11.62 2.125 11.9 2.685 ;
      RECT  12.74 2.125 13.02 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.87 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.87 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.84 -0.14 22.57 0.14 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.91 1.565 13.555 1.795 ;
      RECT  13.325 1.795 13.555 3.805 ;
      RECT  5.43 3.805 16.97 4.035 ;
    END
    ANTENNADIFFAREA 12.316 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.55 0.445 21.45 0.675 ;
      RECT  8.55 0.675 8.78 1.005 ;
      RECT  0.18 1.005 8.78 1.235 ;
      RECT  9.14 1.005 22.22 1.235 ;
      RECT  0.18 4.365 6.835 4.595 ;
      RECT  6.605 4.595 6.835 4.925 ;
      RECT  6.605 4.925 8.01 5.155 ;
      RECT  15.86 4.365 22.22 4.595 ;
      RECT  15.86 4.595 16.09 4.925 ;
      RECT  14.39 4.925 16.09 5.155 ;
  END
END MDN_OAI221_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI22_1
#      Description : Two 2-input ORs into 2-input NAND
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI22_1
  CLASS CORE ;
  FOREIGN MDN_OAI22_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 4.65 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  0.0 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 4.65 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 3.805 ;
      RECT  1.72 3.805 2.76 4.035 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 2.355 0.675 ;
      RECT  2.125 0.675 2.355 1.005 ;
      RECT  2.125 1.005 4.3 1.235 ;
  END
END MDN_OAI22_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI22_2
#      Description : Two 2-input ORs into 2-input NAND
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI22_2
  CLASS CORE ;
  FOREIGN MDN_OAI22_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 4.365 8.78 4.595 ;
      RECT  8.285 4.595 8.515 5.46 ;
      RECT  8.285 5.46 9.13 5.74 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  7.725 0.14 7.955 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 4.035 1.235 ;
      RECT  3.805 1.235 4.035 1.565 ;
      RECT  3.805 1.565 4.595 1.795 ;
      RECT  4.365 1.795 4.595 4.365 ;
      RECT  2.42 4.365 6.54 4.595 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 4.595 0.675 ;
      RECT  4.365 0.675 4.595 1.005 ;
      RECT  4.365 1.005 8.78 1.235 ;
      RECT  0.95 4.925 3.53 5.155 ;
      RECT  5.43 4.925 8.01 5.155 ;
  END
END MDN_OAI22_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI22_3
#      Description : Two 2-input ORs into 2-input NAND
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI22_3
  CLASS CORE ;
  FOREIGN MDN_OAI22_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 6.3 2.355 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 9.66 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 13.02 2.355 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.68 4.365 13.26 4.595 ;
      RECT  12.765 4.595 12.995 5.46 ;
      RECT  12.32 5.46 13.61 5.74 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 6.275 1.235 ;
      RECT  6.045 1.235 6.275 1.565 ;
      RECT  6.045 1.565 6.835 1.795 ;
      RECT  6.605 1.795 6.835 4.365 ;
      RECT  3.96 4.365 9.48 4.595 ;
    END
    ANTENNADIFFAREA 9.072 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 6.835 0.675 ;
      RECT  6.605 0.675 6.835 1.005 ;
      RECT  6.605 1.005 13.26 1.235 ;
      RECT  0.95 4.925 5.77 5.155 ;
      RECT  7.67 4.925 12.49 5.155 ;
  END
END MDN_OAI22_3
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI22_4
#      Description : Two 2-input ORs into 2-input NAND
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI22_4
  CLASS CORE ;
  FOREIGN MDN_OAI22_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.87 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.87 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  8.4 5.46 9.52 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  8.79 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 8.475 1.235 ;
      RECT  8.03 1.235 8.475 1.26 ;
      RECT  8.245 1.26 8.475 1.565 ;
      RECT  8.245 1.565 9.075 1.795 ;
      RECT  8.845 1.795 9.075 4.365 ;
      RECT  4.66 4.365 13.26 4.595 ;
    END
    ANTENNADIFFAREA 12.096 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 9.075 0.675 ;
      RECT  8.845 0.675 9.075 1.005 ;
      RECT  8.845 1.005 17.74 1.235 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  4.07 4.595 4.3 4.925 ;
      RECT  4.07 4.925 8.01 5.155 ;
      RECT  13.62 4.365 17.74 4.595 ;
      RECT  13.62 4.595 13.85 4.925 ;
      RECT  9.91 4.925 13.85 5.155 ;
  END
END MDN_OAI22_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI311_1
#      Description : 3-input OR into 3-input NAND
#      Equation    : X=!((A1|A2|A3)&B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI311_1
  CLASS CORE ;
  FOREIGN MDN_OAI311_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  1.005 5.46 2.41 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      RECT  3.245 0.14 3.475 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 1.005 6.54 1.235 ;
      RECT  5.485 1.235 5.715 3.805 ;
      RECT  3.96 3.805 6.54 4.035 ;
    END
    ANTENNADIFFAREA 3.308 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.005 5.0 1.235 ;
      RECT  1.72 4.365 2.76 4.595 ;
  END
END MDN_OAI311_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI311_2
#      Description : 3-input OR into 3-input NAND
#      Equation    : X=!((A1|A2|A3)&B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI311_2
  CLASS CORE ;
  FOREIGN MDN_OAI311_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.685 ;
      RECT  4.9 2.685 6.3 2.915 ;
      RECT  6.02 2.125 6.3 2.685 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.685 ;
      RECT  9.38 2.685 10.78 2.915 ;
      RECT  10.5 2.125 10.78 2.685 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 7.42 2.685 ;
      RECT  7.14 2.685 8.54 2.915 ;
      RECT  8.26 2.125 8.54 2.685 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.08 -0.14 11.37 0.14 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.405 1.005 11.02 1.235 ;
      RECT  9.405 1.235 9.635 1.565 ;
      RECT  8.845 1.565 9.635 1.795 ;
      RECT  8.845 1.795 9.075 3.805 ;
      RECT  4.66 3.805 11.02 4.035 ;
    END
    ANTENNADIFFAREA 6.616 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  7.67 0.445 10.25 0.675 ;
      RECT  0.18 1.005 8.78 1.235 ;
      RECT  0.18 3.805 4.3 4.035 ;
      RECT  3.19 4.925 5.77 5.155 ;
  END
END MDN_OAI311_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI311_4
#      Description : 3-input OR into 3-input NAND
#      Equation    : X=!((A1|A2|A3)&B1&B2)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI311_4
  CLASS CORE ;
  FOREIGN MDN_OAI311_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.685 ;
      RECT  9.38 2.685 13.02 2.915 ;
      RECT  10.5 2.125 10.78 2.685 ;
      RECT  11.62 2.125 11.9 2.685 ;
      RECT  12.74 2.125 13.02 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.34 2.125 18.62 2.685 ;
      RECT  18.34 2.685 21.98 2.915 ;
      RECT  19.46 2.125 19.74 2.685 ;
      RECT  20.58 2.125 20.86 2.685 ;
      RECT  21.7 2.125 21.98 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 14.14 2.685 ;
      RECT  13.86 2.685 17.5 2.915 ;
      RECT  14.98 2.125 15.26 2.685 ;
      RECT  16.1 2.125 16.38 2.685 ;
      RECT  17.22 2.125 17.5 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 19.155 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 4.65 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  18.07 5.47 18.33 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.84 -0.14 22.57 0.14 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  7.725 -0.14 10.195 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.365 1.005 22.22 1.235 ;
      RECT  18.365 1.235 18.595 1.565 ;
      RECT  17.805 1.565 18.595 1.795 ;
      RECT  17.805 1.795 18.035 3.805 ;
      RECT  9.14 3.805 22.22 4.035 ;
    END
    ANTENNADIFFAREA 13.232 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  14.39 0.445 21.45 0.675 ;
      RECT  0.18 1.005 17.74 1.235 ;
      RECT  15.86 1.235 16.2 1.245 ;
      RECT  0.18 3.805 8.78 4.035 ;
      RECT  5.43 4.925 12.49 5.155 ;
  END
END MDN_OAI311_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI31_1
#      Description : 3-input OR into 2-input NAND
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI31_1
  CLASS CORE ;
  FOREIGN MDN_OAI31_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 4.65 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 2.76 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 1.005 4.3 1.235 ;
      RECT  3.245 1.235 3.475 3.53 ;
    END
    ANTENNADIFFAREA 2.086 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 3.53 0.675 ;
      RECT  1.72 4.365 2.76 4.595 ;
  END
END MDN_OAI31_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI31_2
#      Description : 3-input OR into 2-input NAND
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI31_2
  CLASS CORE ;
  FOREIGN MDN_OAI31_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.685 ;
      RECT  4.9 2.685 6.3 2.915 ;
      RECT  6.02 2.125 6.3 2.685 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 7.42 2.685 ;
      RECT  7.14 2.685 8.54 2.915 ;
      RECT  8.26 2.125 8.54 2.685 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  1.005 5.46 2.41 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 6.89 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      RECT  3.245 0.14 3.475 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.165 1.005 8.78 1.235 ;
      RECT  7.165 1.235 7.395 1.565 ;
      RECT  6.605 1.565 7.395 1.795 ;
      RECT  6.605 1.795 6.835 3.805 ;
      RECT  4.66 3.805 8.78 4.035 ;
    END
    ANTENNADIFFAREA 4.82 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  6.605 0.445 8.01 0.675 ;
      RECT  6.605 0.675 6.835 1.005 ;
      RECT  0.18 1.005 6.835 1.235 ;
      RECT  0.18 3.805 4.3 4.035 ;
      RECT  3.19 4.925 5.77 5.155 ;
  END
END MDN_OAI31_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI31_3
#      Description : 3-input OR into 2-input NAND
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI31_3
  CLASS CORE ;
  FOREIGN MDN_OAI31_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 7.42 2.685 ;
      RECT  7.14 2.685 9.66 2.915 ;
      RECT  8.26 2.125 8.54 2.685 ;
      RECT  9.38 2.125 9.66 2.685 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 6.3 2.355 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 2.125 11.9 2.685 ;
      RECT  11.62 2.685 13.02 2.915 ;
      RECT  12.74 2.125 13.02 2.685 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.765 4.365 13.26 4.595 ;
      RECT  12.765 4.595 12.995 5.46 ;
      RECT  12.765 5.46 13.61 5.74 ;
      RECT  9.965 4.365 11.72 4.595 ;
      RECT  9.965 4.595 10.195 5.46 ;
      RECT  9.965 5.46 11.76 5.74 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.88 -0.14 13.61 0.14 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  8.84 0.14 9.07 1.005 ;
      RECT  8.84 1.005 9.48 1.235 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.525 1.005 13.26 1.235 ;
      RECT  10.525 1.235 10.755 3.245 ;
      RECT  7.67 3.245 12.49 3.475 ;
    END
    ANTENNADIFFAREA 6.258 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  9.965 0.445 12.49 0.675 ;
      RECT  9.965 0.675 10.195 1.565 ;
      RECT  0.18 1.005 8.515 1.235 ;
      RECT  8.285 1.235 8.515 1.565 ;
      RECT  8.285 1.565 10.195 1.795 ;
      RECT  3.96 4.365 9.48 4.595 ;
      RECT  0.95 4.925 5.77 5.155 ;
      RECT  10.47 5.0 11.93 5.23 ;
  END
END MDN_OAI31_3
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI31_4
#      Description : 3-input OR into 2-input NAND
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI31_4
  CLASS CORE ;
  FOREIGN MDN_OAI31_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 9.66 2.685 ;
      RECT  9.38 2.685 13.02 2.915 ;
      RECT  10.5 2.125 10.78 2.685 ;
      RECT  11.62 2.125 11.9 2.685 ;
      RECT  12.74 2.125 13.02 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 14.14 2.685 ;
      RECT  13.86 2.685 17.5 2.915 ;
      RECT  14.98 2.125 15.26 2.685 ;
      RECT  16.1 2.125 16.38 2.685 ;
      RECT  17.22 2.125 17.5 2.685 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 4.905 16.915 5.46 ;
      RECT  16.685 5.46 18.09 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.445 5.46 15.12 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  3.245 5.46 4.65 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.8 -0.14 18.09 0.14 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  7.725 -0.14 10.195 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.445 1.005 17.74 1.235 ;
      RECT  14.445 1.235 14.675 1.565 ;
      RECT  13.325 1.565 14.675 1.795 ;
      RECT  13.325 1.795 13.555 3.805 ;
      RECT  9.14 3.805 17.74 4.035 ;
    END
    ANTENNADIFFAREA 9.64 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  13.325 0.445 16.97 0.675 ;
      RECT  13.325 0.675 13.555 1.005 ;
      RECT  0.18 1.005 13.555 1.235 ;
      RECT  0.18 3.805 8.78 4.035 ;
      RECT  5.43 4.925 12.49 5.155 ;
  END
END MDN_OAI31_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI32_1
#      Description : 3-input OR and 2-input OR into 2-input NAND
#      Equation    : X=!((A1|A2|A3)&(B1|B2))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI32_1
  CLASS CORE ;
  FOREIGN MDN_OAI32_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  4.31 5.46 5.715 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  0.0 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  3.245 0.14 3.475 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 3.805 ;
      RECT  1.72 3.805 2.76 4.035 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 2.355 0.675 ;
      RECT  2.125 0.675 2.355 1.005 ;
      RECT  2.125 1.005 5.0 1.235 ;
      RECT  3.96 4.365 5.0 4.595 ;
  END
END MDN_OAI32_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI32_2
#      Description : 3-input OR and 2-input OR into 2-input NAND
#      Equation    : X=!((A1|A2|A3)&(B1|B2))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI32_2
  CLASS CORE ;
  FOREIGN MDN_OAI32_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 10.78 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 -0.14 11.37 0.14 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.165 1.005 11.02 1.235 ;
      RECT  7.165 1.235 7.395 1.565 ;
      RECT  6.605 1.565 7.395 1.795 ;
      RECT  6.605 1.795 6.835 3.805 ;
      RECT  4.66 3.805 8.78 4.035 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  6.605 0.445 10.25 0.675 ;
      RECT  6.605 0.675 6.835 1.005 ;
      RECT  0.18 1.005 6.835 1.235 ;
      RECT  0.175 4.365 4.3 4.595 ;
      RECT  8.845 4.365 11.02 4.595 ;
      RECT  8.845 4.595 9.075 4.925 ;
      RECT  7.67 4.925 9.075 5.155 ;
      RECT  3.19 4.925 5.77 5.155 ;
  END
END MDN_OAI32_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI32_4
#      Description : 3-input OR and 2-input OR into 2-input NAND
#      Equation    : X=!((A1|A2|A3)&(B1|B2))
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI32_4
  CLASS CORE ;
  FOREIGN MDN_OAI32_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.34 2.125 21.98 2.355 ;
      RECT  18.34 2.355 18.62 2.915 ;
      RECT  19.46 2.355 19.74 2.915 ;
      RECT  20.58 2.355 20.86 2.915 ;
      RECT  21.7 2.355 21.98 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.865 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.87 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  8.79 5.46 9.52 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.84 -0.14 22.57 0.14 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.62 1.005 22.22 1.235 ;
      RECT  17.805 1.235 18.035 3.805 ;
      RECT  17.245 3.805 18.035 4.035 ;
      RECT  17.245 4.035 17.475 4.365 ;
      RECT  9.14 4.365 17.475 4.595 ;
    END
    ANTENNADIFFAREA 12.096 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  13.03 0.445 21.45 0.675 ;
      RECT  13.03 0.675 13.26 1.005 ;
      RECT  0.18 1.005 13.26 1.235 ;
      RECT  0.18 4.365 8.78 4.595 ;
      RECT  18.1 4.365 22.22 4.595 ;
      RECT  18.1 4.595 18.33 4.925 ;
      RECT  14.39 4.925 18.33 5.155 ;
      RECT  5.43 4.925 12.49 5.155 ;
  END
END MDN_OAI32_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI41_1
#      Description : 4-input OR into 2-input NAND
#      Equation    : X=!((A1|A2|A3|A4)&B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI41_1
  CLASS CORE ;
  FOREIGN MDN_OAI41_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A4
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 4.365 6.54 4.595 ;
      RECT  6.045 4.595 6.275 5.46 ;
      RECT  6.045 5.46 6.72 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  1.005 5.46 2.41 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.6 -0.14 6.275 0.14 ;
      RECT  6.045 0.14 6.275 1.005 ;
      RECT  4.66 1.005 6.275 1.235 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      RECT  3.245 0.14 3.475 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 1.565 6.545 1.795 ;
      RECT  5.485 1.795 5.715 3.53 ;
    END
    ANTENNADIFFAREA 2.086 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  4.07 0.445 5.77 0.675 ;
      RECT  4.07 0.675 4.3 1.005 ;
      RECT  1.72 1.005 4.3 1.235 ;
      RECT  1.72 4.365 2.76 4.595 ;
      RECT  3.96 4.365 5.0 4.595 ;
  END
END MDN_OAI41_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI41_2
#      Description : 4-input OR into 2-input NAND
#      Equation    : X=!((A1|A2|A3|A4)&B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI41_2
  CLASS CORE ;
  FOREIGN MDN_OAI41_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A4
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 10.78 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.64 -0.14 11.37 0.14 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.845 1.565 10.25 1.795 ;
      RECT  8.845 1.795 9.075 4.365 ;
      RECT  6.9 4.365 11.02 4.595 ;
    END
    ANTENNADIFFAREA 4.686 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 11.02 1.235 ;
      RECT  2.42 4.365 6.54 4.595 ;
      RECT  0.95 4.925 3.53 5.155 ;
      RECT  5.43 4.925 8.01 5.155 ;
  END
END MDN_OAI41_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OAI41_4
#      Description : 4-input OR into 2-input NAND
#      Equation    : X=!((A1|A2|A3|A4)&B)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAI41_4
  CLASS CORE ;
  FOREIGN MDN_OAI41_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.065 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A4
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.34 2.125 21.98 2.355 ;
      RECT  18.34 2.355 18.62 2.915 ;
      RECT  19.46 2.355 19.74 2.915 ;
      RECT  20.58 2.355 20.86 2.915 ;
      RECT  21.7 2.355 21.98 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  10.64 5.46 11.76 5.74 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.84 -0.14 22.57 0.14 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.73 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.73 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  10.64 -0.14 11.76 0.14 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  18.365 1.005 22.22 1.235 ;
      RECT  18.365 1.235 18.595 1.565 ;
      RECT  17.805 1.565 18.595 1.795 ;
      RECT  17.805 1.795 18.035 4.365 ;
      RECT  13.62 4.365 22.22 4.595 ;
    END
    ANTENNADIFFAREA 9.64 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  17.805 0.445 21.45 0.675 ;
      RECT  17.805 0.675 18.035 1.005 ;
      RECT  0.14 1.005 18.035 1.235 ;
      RECT  0.18 4.365 8.78 4.595 ;
      RECT  9.1 4.365 13.26 4.595 ;
      RECT  13.03 4.595 13.26 4.925 ;
      RECT  13.03 4.925 16.97 5.155 ;
      RECT  5.43 4.925 12.49 5.155 ;
  END
END MDN_OAI41_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OAOI211_1
#      Description : One 2-input OR into 2-input AND into 2-input NOR
#      Equation    : X=!(((A1|A2)&B)|C)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAOI211_1
  CLASS CORE ;
  FOREIGN MDN_OAOI211_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.36 5.46 4.035 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 1.12 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 2.76 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 1.51 3.475 4.365 ;
      RECT  2.42 4.365 3.475 4.595 ;
    END
    ANTENNADIFFAREA 1.992 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.95 0.445 4.035 0.675 ;
      RECT  3.805 0.675 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  1.72 4.365 2.06 4.595 ;
      RECT  1.83 4.595 2.06 4.925 ;
      RECT  1.83 4.925 3.53 5.155 ;
  END
END MDN_OAOI211_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OAOI211_2
#      Description : One 2-input OR into 2-input AND into 2-input NOR
#      Equation    : X=!(((A1|A2)&B)|C)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAOI211_2
  CLASS CORE ;
  FOREIGN MDN_OAOI211_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.87 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.005 8.78 1.235 ;
      RECT  6.605 1.235 6.835 3.245 ;
      RECT  6.605 3.245 8.01 3.475 ;
    END
    ANTENNADIFFAREA 3.928 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  4.07 0.445 5.77 0.675 ;
      RECT  4.07 0.675 4.3 1.005 ;
      RECT  0.18 1.005 4.3 1.235 ;
      RECT  8.285 4.365 8.78 4.595 ;
      RECT  8.285 4.595 8.515 4.925 ;
      RECT  2.42 4.365 7.395 4.595 ;
      RECT  7.165 4.595 7.395 4.925 ;
      RECT  7.165 4.925 8.515 5.155 ;
      RECT  0.95 4.925 3.53 5.155 ;
  END
END MDN_OAOI211_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OAOI211_3
#      Description : One 2-input OR into 2-input AND into 2-input NOR
#      Equation    : X=!(((A1|A2)&B)|C)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAOI211_3
  CLASS CORE ;
  FOREIGN MDN_OAOI211_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 6.3 2.355 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 9.66 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 13.02 2.355 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.88 5.46 13.61 5.74 ;
      RECT  9.14 4.365 9.635 4.595 ;
      RECT  9.405 4.595 9.635 5.46 ;
      RECT  7.725 4.87 7.955 5.46 ;
      RECT  7.725 5.46 9.635 5.74 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.32 -0.14 13.61 0.14 ;
      RECT  12.765 0.14 12.995 1.005 ;
      RECT  10.68 1.005 13.26 1.235 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.245 -0.14 3.92 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.67 0.445 12.49 0.675 ;
      RECT  9.965 0.675 10.195 3.245 ;
      RECT  9.965 3.245 10.755 3.475 ;
      RECT  10.525 3.475 10.755 4.365 ;
      RECT  10.525 4.365 13.26 4.595 ;
    END
    ANTENNADIFFAREA 5.976 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 9.48 1.235 ;
      RECT  8.55 3.805 10.195 4.035 ;
      RECT  8.55 4.035 8.78 4.365 ;
      RECT  9.965 4.035 10.195 4.925 ;
      RECT  3.96 4.365 8.78 4.595 ;
      RECT  9.965 4.925 12.49 5.155 ;
      RECT  0.95 4.925 5.77 5.155 ;
  END
END MDN_OAOI211_3
#-----------------------------------------------------------------------
#      Cell        : MDN_OAOI211_4
#      Description : One 2-input OR into 2-input AND into 2-input NOR
#      Equation    : X=!(((A1|A2)&B)|C)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OAOI211_4
  CLASS CORE ;
  FOREIGN MDN_OAOI211_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.92 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 8.54 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 4.06 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  13.86 2.125 17.5 2.355 ;
      RECT  13.86 2.355 14.14 2.915 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
      RECT  17.22 2.355 17.5 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  17.36 5.46 18.09 5.74 ;
      RECT  9.965 4.87 10.195 5.46 ;
      RECT  9.965 5.46 12.435 5.74 ;
      RECT  12.205 4.87 12.435 5.46 ;
      RECT  3.245 4.87 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 17.92 5.74 ;
      LAYER VIA12 ;
      RECT  17.51 5.47 17.77 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  16.685 -0.14 18.09 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.445 -0.14 15.12 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  7.725 -0.14 8.4 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 17.92 0.14 ;
      LAYER VIA12 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  17.51 -0.13 17.77 0.13 ;
      RECT  14.71 -0.13 14.97 0.13 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.14 1.005 17.74 1.235 ;
      RECT  13.325 1.235 13.555 3.245 ;
      RECT  13.325 3.245 16.97 3.475 ;
    END
    ANTENNADIFFAREA 8.18 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.55 0.445 12.49 0.675 ;
      RECT  8.55 0.675 8.78 1.005 ;
      RECT  0.18 1.005 8.78 1.235 ;
      RECT  0.18 4.365 8.78 4.595 ;
      RECT  15.565 4.365 17.74 4.595 ;
      RECT  15.565 4.595 15.795 4.925 ;
      RECT  9.14 4.365 13.555 4.595 ;
      RECT  9.14 4.595 9.37 4.925 ;
      RECT  13.325 4.595 13.555 4.925 ;
      RECT  5.43 4.925 9.37 5.155 ;
      RECT  13.325 4.925 15.795 5.155 ;
  END
END MDN_OAOI211_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OR2_1
#      Description : 2-Input OR
#      Equation    : X=A1|A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR2_1
  CLASS CORE ;
  FOREIGN MDN_OR2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      RECT  3.245 0.14 3.475 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.09 0.6 ;
      RECT  3.75 0.6 3.98 1.005 ;
      RECT  0.18 1.005 3.98 1.235 ;
      RECT  2.125 1.235 2.355 3.245 ;
      RECT  1.72 3.245 2.355 3.475 ;
  END
END MDN_OR2_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OR2_12
#      Description : 2-Input OR
#      Equation    : X=A1|A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR2_12
  CLASS CORE ;
  FOREIGN MDN_OR2_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 6.3 2.355 ;
      RECT  3.78 2.355 4.06 2.915 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 2.94 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
      RECT  2.66 2.355 2.94 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 20.33 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.24 5.46 16.915 5.74 ;
      RECT  14.445 4.9 14.675 5.46 ;
      RECT  14.0 5.46 14.675 5.74 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 12.88 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  6.55 5.46 7.955 5.74 ;
      RECT  0.18 4.365 2.76 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 1.12 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 20.16 5.74 ;
      LAYER VIA12 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  19.75 5.47 20.01 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  14.15 5.47 14.41 5.73 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  18.925 -0.14 20.33 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.685 -0.14 17.36 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  14.0 -0.14 14.675 0.14 ;
      RECT  14.445 0.14 14.675 0.7 ;
      RECT  12.205 -0.14 12.88 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 20.16 0.14 ;
      LAYER VIA12 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  19.75 -0.13 20.01 0.13 ;
      RECT  16.95 -0.13 17.21 0.13 ;
      RECT  14.15 -0.13 14.41 0.13 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.955 1.4 19.925 1.96 ;
      RECT  17.64 1.96 18.2 3.08 ;
      RECT  6.955 3.08 19.925 3.64 ;
    END
    ANTENNADIFFAREA 18.144 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  6.31 0.37 7.45 0.6 ;
      RECT  6.31 0.6 6.54 1.005 ;
      RECT  0.18 1.005 6.54 1.235 ;
      RECT  17.19 0.37 18.65 0.6 ;
      RECT  7.11 2.405 17.41 2.635 ;
      RECT  18.43 2.405 19.77 2.635 ;
      RECT  3.96 4.365 6.835 4.595 ;
      RECT  6.605 4.595 6.835 5.0 ;
      RECT  6.605 5.0 7.45 5.23 ;
      RECT  0.95 4.925 5.77 5.155 ;
  END
END MDN_OR2_12
#-----------------------------------------------------------------------
#      Cell        : MDN_OR2_2
#      Description : 2-Input OR
#      Equation    : X=A1|A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR2_2
  CLASS CORE ;
  FOREIGN MDN_OR2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      RECT  3.245 0.14 3.475 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 4.3 1.795 ;
      RECT  3.245 1.795 3.475 3.245 ;
      RECT  2.42 3.245 4.3 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.09 0.6 ;
      RECT  3.75 0.6 3.98 1.005 ;
      RECT  2.63 0.37 2.97 0.6 ;
      RECT  2.63 0.6 2.86 1.005 ;
      RECT  0.18 1.005 3.98 1.235 ;
      RECT  1.565 1.235 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
  END
END MDN_OR2_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OR2_3
#      Description : 2-Input OR
#      Equation    : X=A1|A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR2_3
  CLASS CORE ;
  FOREIGN MDN_OR2_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  3.245 0.14 3.475 0.7 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.565 5.0 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  2.42 3.245 5.0 3.475 ;
    END
    ANTENNADIFFAREA 4.536 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 5.21 0.6 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.405 ;
      RECT  1.565 2.405 4.09 2.635 ;
      RECT  1.565 2.635 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
  END
END MDN_OR2_3
#-----------------------------------------------------------------------
#      Cell        : MDN_OR2_4
#      Description : 2-Input OR
#      Equation    : X=A1|A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR2_4
  CLASS CORE ;
  FOREIGN MDN_OR2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 5.715 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      RECT  3.245 0.14 3.475 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 2.915 1.235 ;
      RECT  2.685 1.235 2.915 1.565 ;
      RECT  2.685 1.565 6.54 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  2.685 3.245 6.54 3.475 ;
      RECT  2.685 3.475 2.915 3.805 ;
      RECT  2.42 3.805 2.915 4.035 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.98 0.6 5.21 1.005 ;
      RECT  4.98 1.005 6.22 1.235 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 2.405 ;
      RECT  2.125 2.405 5.04 2.635 ;
      RECT  2.125 2.635 2.355 3.245 ;
      RECT  1.72 3.245 2.355 3.475 ;
  END
END MDN_OR2_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OR2_6
#      Description : 2-Input OR
#      Equation    : X=A1|A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR2_6
  CLASS CORE ;
  FOREIGN MDN_OR2_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 11.37 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  9.11 -0.13 9.37 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 0.98 5.735 1.26 ;
      RECT  5.455 1.26 5.735 1.54 ;
      RECT  5.455 1.54 11.02 1.82 ;
      RECT  8.82 1.82 9.1 3.22 ;
      RECT  5.46 3.22 11.02 3.5 ;
      RECT  5.46 3.5 5.74 4.34 ;
      RECT  4.66 4.34 5.74 4.62 ;
    END
    ANTENNADIFFAREA 9.072 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  8.23 0.37 9.69 0.6 ;
      RECT  0.18 1.005 4.035 1.235 ;
      RECT  3.805 1.235 4.035 1.565 ;
      RECT  3.805 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 2.405 ;
      RECT  4.925 2.405 8.57 2.635 ;
      RECT  4.925 2.635 5.155 3.805 ;
      RECT  3.805 3.805 5.155 4.035 ;
      RECT  3.805 4.035 4.035 4.365 ;
      RECT  2.42 4.365 4.035 4.595 ;
      RECT  9.35 2.405 10.81 2.635 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  1.83 4.595 2.06 4.925 ;
      RECT  1.83 4.925 3.53 5.155 ;
  END
END MDN_OR2_6
#-----------------------------------------------------------------------
#      Cell        : MDN_OR2_8
#      Description : 2-Input OR
#      Equation    : X=A1|A2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR2_8
  CLASS CORE ;
  FOREIGN MDN_OR2_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.52 5.46 10.195 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.715 1.495 13.205 1.865 ;
      RECT  11.015 1.865 11.385 3.175 ;
      RECT  4.715 3.175 13.205 3.545 ;
    END
    ANTENNADIFFAREA 12.096 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  4.365 0.37 5.21 0.6 ;
      RECT  4.365 0.6 4.595 1.005 ;
      RECT  0.18 1.005 4.595 1.235 ;
      RECT  4.87 2.405 10.785 2.635 ;
      RECT  11.615 2.405 13.05 2.635 ;
      RECT  0.18 4.365 2.06 4.595 ;
      RECT  1.83 4.595 2.06 4.925 ;
      RECT  1.83 4.925 3.53 5.155 ;
      RECT  2.42 4.365 4.595 4.595 ;
      RECT  4.365 4.595 4.595 5.0 ;
      RECT  4.365 5.0 5.21 5.23 ;
      RECT  10.47 5.0 11.93 5.23 ;
  END
END MDN_OR2_8
#-----------------------------------------------------------------------
#      Cell        : MDN_OR3_1
#      Description : 3-Input OR
#      Equation    : X=A1|A2|A3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR3_1
  CLASS CORE ;
  FOREIGN MDN_OR3_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 4.365 0.7 5.0 ;
      RECT  0.39 5.0 0.73 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.07 5.46 3.475 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 4.65 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  0.56 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  3.75 0.37 4.09 0.6 ;
      RECT  3.75 0.6 3.98 1.005 ;
      RECT  0.18 1.005 3.98 1.235 ;
      RECT  0.445 1.235 0.675 3.245 ;
      RECT  0.18 3.245 0.675 3.475 ;
      RECT  1.72 4.365 2.765 4.595 ;
  END
END MDN_OR3_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OR3_2
#      Description : 3-Input OR
#      Equation    : X=A1|A2|A3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR3_2
  CLASS CORE ;
  FOREIGN MDN_OR3_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 4.365 4.06 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  1.005 5.46 2.8 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.245 0.14 3.475 0.735 ;
      RECT  1.005 -0.14 1.68 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 6.54 1.795 ;
      RECT  5.485 1.795 5.715 3.245 ;
      RECT  4.66 3.245 6.54 3.475 ;
    END
    ANTENNADIFFAREA 3.024 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  5.99 0.6 6.22 1.005 ;
      RECT  4.87 0.37 5.21 0.6 ;
      RECT  4.87 0.6 5.1 1.005 ;
      RECT  1.72 1.005 6.22 1.235 ;
      RECT  3.805 1.235 4.035 3.245 ;
      RECT  3.805 3.245 4.305 3.475 ;
      RECT  1.72 4.365 2.76 4.595 ;
  END
END MDN_OR3_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OR3_4
#      Description : 3-Input OR
#      Equation    : X=A1|A2|A3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR3_4
  CLASS CORE ;
  FOREIGN MDN_OR3_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 4.365 4.06 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.91 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 7.955 0.14 ;
      RECT  5.485 0.14 5.715 0.7 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  1.005 -0.14 1.68 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  6.87 -0.13 7.13 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.565 8.785 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  4.66 3.245 8.78 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 7.45 0.6 ;
      RECT  1.72 1.005 4.3 1.235 ;
      RECT  3.805 1.235 4.035 2.39 ;
      RECT  3.805 2.39 6.145 2.62 ;
      RECT  3.805 2.62 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
      RECT  7.11 2.39 8.42 2.62 ;
      RECT  1.72 4.365 2.77 4.595 ;
  END
END MDN_OR3_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OR3_6
#      Description : 3-Input OR
#      Equation    : X=A1|A2|A3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR3_6
  CLASS CORE ;
  FOREIGN MDN_OR3_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 4.06 2.355 ;
      RECT  2.66 2.355 2.94 2.915 ;
      RECT  3.78 2.355 4.06 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 1.82 2.355 ;
      RECT  0.42 2.355 0.7 2.915 ;
      RECT  1.54 2.355 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.7 ;
      RECT  9.52 -0.14 10.195 0.14 ;
      RECT  9.965 0.14 10.195 0.7 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.7 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  9.67 -0.13 9.93 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.9 1.005 7.42 1.235 ;
      RECT  7.14 1.235 7.42 1.54 ;
      RECT  7.14 1.54 13.26 1.82 ;
      RECT  11.06 1.82 11.34 3.22 ;
      RECT  7.14 3.22 13.26 3.5 ;
      RECT  7.14 3.5 7.42 3.805 ;
      RECT  6.9 3.805 7.42 4.035 ;
    END
    ANTENNADIFFAREA 9.072 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.175 1.005 6.275 1.235 ;
      RECT  6.045 1.235 6.275 1.565 ;
      RECT  6.045 1.565 6.835 1.795 ;
      RECT  6.605 1.795 6.835 2.39 ;
      RECT  6.605 2.39 10.81 2.62 ;
      RECT  6.605 2.62 6.835 3.245 ;
      RECT  6.005 3.245 6.835 3.475 ;
      RECT  6.005 3.475 6.235 3.805 ;
      RECT  4.66 3.805 6.235 4.035 ;
      RECT  11.59 2.39 13.05 2.62 ;
      RECT  0.18 3.805 4.3 4.035 ;
      RECT  3.19 4.925 5.77 5.155 ;
      RECT  10.47 5.0 11.94 5.23 ;
  END
END MDN_OR3_6
#-----------------------------------------------------------------------
#      Cell        : MDN_OR3B_1
#      Description : 3-Input OR (A inverted input)
#      Equation    : X=!A|B1|B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR3B_1
  CLASS CORE ;
  FOREIGN MDN_OR3B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 4.365 4.3 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 4.65 5.74 ;
      RECT  2.42 4.365 2.915 4.595 ;
      RECT  2.685 4.595 2.915 5.46 ;
      RECT  2.24 5.46 2.915 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  0.0 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  3.805 -0.14 4.65 0.14 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  1.005 -0.14 1.68 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.42 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 3.53 ;
    END
    ANTENNADIFFAREA 2.086 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
  END
END MDN_OR3B_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OR3B_2
#      Description : 3-Input OR (A inverted input)
#      Equation    : X=!A|B1|B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR3B_2
  CLASS CORE ;
  FOREIGN MDN_OR3B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 6.3 2.355 ;
      RECT  4.9 2.355 5.18 2.915 ;
      RECT  6.02 2.355 6.3 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  2.8 5.46 3.475 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  1.005 -0.14 2.41 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 1.51 3.475 3.805 ;
      RECT  2.42 3.805 4.595 4.035 ;
      RECT  4.365 4.035 4.595 4.365 ;
      RECT  4.365 4.365 6.54 4.595 ;
    END
    ANTENNADIFFAREA 4.686 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.565 0.37 4.09 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.92 1.795 ;
      RECT  2.69 1.795 2.92 3.245 ;
      RECT  1.72 3.245 2.92 3.475 ;
      RECT  2.42 1.005 6.54 1.235 ;
  END
END MDN_OR3B_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OR3B_3
#      Description : 3-Input OR (A inverted input)
#      Equation    : X=!A|B1|B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR3B_3
  CLASS CORE ;
  FOREIGN MDN_OR3B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 8.54 2.355 ;
      RECT  6.02 2.355 6.3 2.915 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.84 -0.14 9.13 0.14 ;
      RECT  8.285 0.14 8.515 1.005 ;
      RECT  6.2 1.005 8.78 1.235 ;
      RECT  1.005 -0.14 1.68 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.19 1.565 5.0 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  2.42 3.245 4.595 3.475 ;
      RECT  4.365 3.475 4.595 3.805 ;
      RECT  4.365 3.805 8.78 4.035 ;
    END
    ANTENNADIFFAREA 7.096 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.565 0.37 5.21 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  5.485 0.445 8.01 0.675 ;
      RECT  5.485 0.675 5.715 1.005 ;
      RECT  2.42 1.005 5.715 1.235 ;
  END
END MDN_OR3B_3
#-----------------------------------------------------------------------
#      Cell        : MDN_OR3B_4
#      Description : 3-Input OR (A inverted input)
#      Equation    : X=!A|B1|B2
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR3B_4
  CLASS CORE ;
  FOREIGN MDN_OR3B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 10.78 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.725 5.46 8.4 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.99 5.47 8.25 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  7.28 -0.14 7.955 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  7.43 -0.13 7.69 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.19 1.565 5.77 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  2.42 3.245 6.835 3.475 ;
      RECT  6.605 3.475 6.835 3.805 ;
      RECT  6.605 3.805 11.02 4.035 ;
    END
    ANTENNADIFFAREA 9.372 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.565 0.37 6.33 0.6 ;
      RECT  1.565 0.6 1.795 1.005 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  2.42 1.005 11.02 1.235 ;
  END
END MDN_OR3B_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OR4_1
#      Description : 4-Input OR
#      Equation    : X=A1|A2|A3|A4
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR4_1
  CLASS CORE ;
  FOREIGN MDN_OR4_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 4.365 5.18 5.0 ;
      RECT  4.87 5.0 5.21 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 4.365 1.82 5.0 ;
      RECT  1.51 5.0 1.85 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 4.365 6.54 4.595 ;
      RECT  6.045 4.595 6.275 5.46 ;
      RECT  6.045 5.46 6.89 5.74 ;
      RECT  3.245 4.9 3.475 5.46 ;
      RECT  3.245 5.46 3.92 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  3.51 5.47 3.77 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  5.485 -0.14 6.89 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  -0.17 -0.14 2.41 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      RECT  2.125 0.14 2.355 1.005 ;
      RECT  2.125 1.005 2.76 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.245 1.565 4.3 1.795 ;
      RECT  3.245 1.795 3.475 3.245 ;
      RECT  2.42 3.245 4.3 3.475 ;
    END
    ANTENNADIFFAREA 2.41 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.06 1.795 ;
      RECT  1.565 1.795 1.795 2.39 ;
      RECT  1.565 2.39 2.785 2.62 ;
      RECT  1.565 2.62 1.795 3.245 ;
      RECT  1.565 3.245 2.06 3.475 ;
      RECT  4.925 1.005 6.54 1.235 ;
      RECT  4.925 1.235 5.155 1.565 ;
      RECT  4.66 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 2.685 ;
      RECT  3.805 2.39 4.035 2.685 ;
      RECT  3.805 2.685 5.155 2.915 ;
      RECT  4.925 2.915 5.155 3.245 ;
      RECT  4.66 3.245 5.155 3.475 ;
  END
END MDN_OR4_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OR4_2
#      Description : 4-Input OR
#      Equation    : X=A1|A2|A3|A4
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR4_2
  CLASS CORE ;
  FOREIGN MDN_OR4_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 7.42 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.26 2.125 8.54 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  8.285 4.365 8.78 4.595 ;
      RECT  8.285 4.595 8.515 5.46 ;
      RECT  8.285 5.46 9.13 5.74 ;
      RECT  6.045 4.365 6.54 4.595 ;
      RECT  6.045 4.595 6.275 5.46 ;
      RECT  6.045 5.46 6.72 5.74 ;
      RECT  3.805 4.365 5.0 4.595 ;
      RECT  3.805 4.595 4.035 5.46 ;
      RECT  3.805 5.46 4.65 5.74 ;
      RECT  2.42 4.365 2.915 4.595 ;
      RECT  2.685 4.595 2.915 5.46 ;
      RECT  2.24 5.46 2.915 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  1.005 -0.14 1.68 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.365 1.565 5.72 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  3.19 3.245 5.795 3.475 ;
    END
    ANTENNADIFFAREA 4.038 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 1.755 1.235 ;
      RECT  1.525 1.235 1.755 1.565 ;
      RECT  1.52 1.565 2.355 1.795 ;
      RECT  2.125 1.795 2.355 2.39 ;
      RECT  2.125 2.39 3.995 2.62 ;
      RECT  2.125 2.62 2.355 3.245 ;
      RECT  1.72 3.245 2.355 3.475 ;
      RECT  2.42 1.005 6.54 1.235 ;
      RECT  7.15 1.005 8.78 1.235 ;
      RECT  7.15 1.235 7.38 1.565 ;
      RECT  6.605 1.565 7.38 1.795 ;
      RECT  6.605 1.795 6.835 2.39 ;
      RECT  4.87 2.39 6.835 2.62 ;
      RECT  6.605 2.62 6.835 3.245 ;
      RECT  6.605 3.245 7.24 3.475 ;
  END
END MDN_OR4_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OR4_4
#      Description : 4-Input OR
#      Equation    : X=A1|A2|A3|A4
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR4_4
  CLASS CORE ;
  FOREIGN MDN_OR4_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  11.62 2.125 11.9 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  12.74 2.125 13.02 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.765 4.365 13.26 4.595 ;
      RECT  12.765 4.595 12.995 5.46 ;
      RECT  12.765 5.46 13.61 5.74 ;
      RECT  10.525 4.365 11.02 4.595 ;
      RECT  10.525 4.595 10.755 5.46 ;
      RECT  10.525 5.46 11.2 5.74 ;
      RECT  8.44 4.365 9.635 4.595 ;
      RECT  9.405 4.595 9.635 5.46 ;
      RECT  8.4 5.46 9.635 5.74 ;
      RECT  6.2 4.365 7.395 4.595 ;
      RECT  7.165 4.595 7.395 5.46 ;
      RECT  6.16 5.46 7.395 5.74 ;
      RECT  3.96 4.365 5.155 4.595 ;
      RECT  4.925 4.595 5.155 5.46 ;
      RECT  3.92 5.46 5.155 5.74 ;
      RECT  2.42 4.365 2.915 4.595 ;
      RECT  2.685 4.595 2.915 5.46 ;
      RECT  2.24 5.46 2.915 5.74 ;
      RECT  0.18 4.365 0.675 4.595 ;
      RECT  0.445 4.595 0.675 5.46 ;
      RECT  -0.17 5.46 0.675 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  9.11 5.47 9.37 5.73 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  4.07 5.47 4.33 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  5.04 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.73 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.605 1.565 10.25 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  3.19 3.245 10.25 3.475 ;
    END
    ANTENNADIFFAREA 8.076 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  0.18 1.005 1.795 1.235 ;
      RECT  1.565 1.235 1.795 1.565 ;
      RECT  1.565 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 2.685 ;
      RECT  2.685 2.685 6.275 2.915 ;
      RECT  3.805 2.33 4.035 2.685 ;
      RECT  4.925 2.335 5.155 2.685 ;
      RECT  6.045 2.335 6.275 2.685 ;
      RECT  2.685 2.915 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
      RECT  2.42 1.005 11.02 1.235 ;
      RECT  11.645 1.005 13.26 1.235 ;
      RECT  11.645 1.235 11.875 1.565 ;
      RECT  10.525 1.565 11.875 1.795 ;
      RECT  10.525 1.795 10.755 2.685 ;
      RECT  7.165 2.335 7.395 2.685 ;
      RECT  7.16 2.685 10.755 2.915 ;
      RECT  8.285 2.335 8.515 2.685 ;
      RECT  9.405 2.335 9.635 2.685 ;
      RECT  10.525 2.915 10.755 3.245 ;
      RECT  10.525 3.245 11.72 3.475 ;
  END
END MDN_OR4_4
#-----------------------------------------------------------------------
#      Cell        : MDN_OR4B_1
#      Description : 4-Input OR (A inverted input)
#      Equation    : X=!A|B1|B2|B3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR4B_1
  CLASS CORE ;
  FOREIGN MDN_OR4B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  6.02 2.125 6.3 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 4.365 6.54 4.595 ;
      RECT  6.045 4.595 6.275 5.46 ;
      RECT  6.045 5.46 6.89 5.74 ;
      RECT  4.66 4.365 5.155 4.595 ;
      RECT  4.925 4.595 5.155 5.46 ;
      RECT  4.48 5.46 5.155 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  1.005 5.46 1.68 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 6.72 5.74 ;
      LAYER VIA12 ;
      RECT  6.31 5.47 6.57 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  6.045 -0.14 6.89 0.14 ;
      RECT  6.045 0.14 6.275 1.005 ;
      RECT  6.045 1.005 6.54 1.235 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  1.005 -0.14 1.68 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 6.72 0.14 ;
      LAYER VIA12 ;
      RECT  6.31 -0.13 6.57 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.005 5.155 1.235 ;
      RECT  4.925 1.235 5.155 3.245 ;
      RECT  4.925 3.245 5.77 3.475 ;
    END
    ANTENNADIFFAREA 2.086 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  4.87 0.37 5.21 0.445 ;
      RECT  4.015 0.445 5.21 0.675 ;
      RECT  4.015 0.675 4.245 1.005 ;
      RECT  1.72 1.005 4.245 1.235 ;
      RECT  4.015 1.235 4.245 1.565 ;
      RECT  4.015 1.565 4.595 1.795 ;
      RECT  4.365 1.795 4.595 3.245 ;
      RECT  3.96 3.245 4.595 3.475 ;
      RECT  1.72 4.365 2.76 4.595 ;
  END
END MDN_OR4B_1
#-----------------------------------------------------------------------
#      Cell        : MDN_OR4B_2
#      Description : 4-Input OR (A inverted input)
#      Equation    : X=!A|B1|B2|B3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR4B_2
  CLASS CORE ;
  FOREIGN MDN_OR4B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.96 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.14 2.125 8.54 2.355 ;
      RECT  7.14 2.355 7.42 2.915 ;
      RECT  8.26 2.355 8.54 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 2.125 4.06 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  8.285 4.365 8.78 4.595 ;
      RECT  8.285 4.595 8.515 5.46 ;
      RECT  8.285 5.46 9.13 5.74 ;
      RECT  6.2 4.365 7.395 4.595 ;
      RECT  7.165 4.595 7.395 5.46 ;
      RECT  6.55 5.46 7.395 5.74 ;
      RECT  4.66 4.365 5.155 4.595 ;
      RECT  4.925 4.595 5.155 5.46 ;
      RECT  4.48 5.46 5.155 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  1.005 5.46 1.68 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 8.96 5.74 ;
      LAYER VIA12 ;
      RECT  8.55 5.47 8.81 5.73 ;
      RECT  6.87 5.47 7.13 5.73 ;
      RECT  4.63 5.47 4.89 5.73 ;
      RECT  1.27 5.47 1.53 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 -0.14 9.13 0.14 ;
      RECT  7.725 0.14 7.955 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  1.005 -0.14 1.68 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 8.96 0.14 ;
      LAYER VIA12 ;
      RECT  7.99 -0.13 8.25 0.13 ;
      RECT  8.55 -0.13 8.81 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  1.27 -0.13 1.53 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.66 1.005 6.275 1.235 ;
      RECT  6.045 1.235 6.275 1.565 ;
      RECT  6.045 1.565 6.835 1.795 ;
      RECT  6.605 1.795 6.835 3.245 ;
      RECT  5.43 3.245 8.01 3.475 ;
    END
    ANTENNADIFFAREA 4.172 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.445 6.835 0.675 ;
      RECT  6.605 0.675 6.835 1.005 ;
      RECT  6.605 1.005 8.78 1.235 ;
      RECT  1.72 1.005 4.3 1.235 ;
      RECT  4.07 1.235 4.3 1.565 ;
      RECT  4.07 1.565 5.155 1.795 ;
      RECT  4.925 1.795 5.155 2.125 ;
      RECT  4.925 2.125 6.275 2.355 ;
      RECT  6.045 2.355 6.275 2.675 ;
      RECT  4.925 2.355 5.155 3.245 ;
      RECT  3.96 3.245 5.155 3.475 ;
      RECT  1.72 4.365 2.76 4.595 ;
  END
END MDN_OR4B_2
#-----------------------------------------------------------------------
#      Cell        : MDN_OR4B_3
#      Description : 4-Input OR (A inverted input)
#      Equation    : X=!A|B1|B2|B3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR4B_3
  CLASS CORE ;
  FOREIGN MDN_OR4B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  8.255 2.125 10.78 2.355 ;
      RECT  8.26 2.355 8.54 2.915 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
    END
    ANTENNAGATEAREA 1.701 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 4.365 4.06 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 11.37 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 11.2 5.74 ;
      LAYER VIA12 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  10.08 -0.14 11.37 0.14 ;
      RECT  10.525 0.14 10.755 1.005 ;
      RECT  8.44 1.005 11.02 1.235 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 11.2 0.14 ;
      LAYER VIA12 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  7.725 1.56 7.955 1.565 ;
      RECT  4.66 1.565 7.955 1.795 ;
      RECT  7.725 1.795 7.955 3.245 ;
      RECT  4.66 3.245 7.96 3.475 ;
      RECT  7.725 3.475 7.955 3.805 ;
      RECT  7.725 3.805 11.02 4.035 ;
    END
    ANTENNADIFFAREA 7.23 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.445 10.25 0.675 ;
      RECT  1.72 1.005 4.035 1.235 ;
      RECT  3.805 1.235 4.035 1.565 ;
      RECT  3.805 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 2.125 ;
      RECT  3.805 2.125 7.395 2.355 ;
      RECT  4.925 2.355 5.155 2.675 ;
      RECT  6.045 2.355 6.275 2.675 ;
      RECT  7.165 2.355 7.395 2.675 ;
      RECT  3.805 2.355 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
      RECT  1.715 4.365 2.76 4.595 ;
  END
END MDN_OR4B_3
#-----------------------------------------------------------------------
#      Cell        : MDN_OR4B_4
#      Description : 4-Input OR (A inverted input)
#      Equation    : X=!A|B1|B2|B3
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_OR4B_4
  CLASS CORE ;
  FOREIGN MDN_OR4B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  9.38 2.125 13.02 2.355 ;
      RECT  9.38 2.355 9.66 2.915 ;
      RECT  10.5 2.355 10.78 2.915 ;
      RECT  11.62 2.355 11.9 2.915 ;
      RECT  12.74 2.355 13.02 2.915 ;
    END
    ANTENNAGATEAREA 2.268 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  3.78 4.365 4.06 5.0 ;
      RECT  3.75 5.0 4.09 5.23 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 4.9 12.435 5.46 ;
      RECT  12.205 5.46 13.61 5.74 ;
      RECT  9.965 4.9 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  7.725 4.9 7.955 5.46 ;
      RECT  7.28 5.46 7.955 5.74 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.9 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 13.44 5.74 ;
      LAYER VIA12 ;
      RECT  12.47 5.47 12.73 5.73 ;
      RECT  13.03 5.47 13.29 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  7.43 5.47 7.69 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  12.205 -0.14 13.61 0.14 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  9.965 -0.14 10.64 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  2.8 -0.14 3.475 0.14 ;
      RECT  3.245 0.14 3.475 0.73 ;
      RECT  -0.17 -0.14 1.235 0.14 ;
      RECT  1.005 0.14 1.235 0.7 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 13.44 0.14 ;
      LAYER VIA12 ;
      RECT  12.47 -0.13 12.73 0.13 ;
      RECT  13.03 -0.13 13.29 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
      RECT  0.71 -0.13 0.97 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.65 1.565 9.075 1.795 ;
      RECT  8.845 1.795 9.075 3.245 ;
      RECT  4.66 3.245 9.075 3.475 ;
      RECT  8.845 3.475 9.075 3.805 ;
      RECT  8.845 3.805 13.26 4.035 ;
    END
    ANTENNADIFFAREA 9.64 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  5.43 0.445 9.33 0.675 ;
      RECT  9.1 0.675 9.33 1.005 ;
      RECT  9.1 1.005 13.26 1.235 ;
      RECT  1.72 1.005 4.035 1.235 ;
      RECT  3.805 1.235 4.035 1.565 ;
      RECT  3.805 1.565 4.3 1.795 ;
      RECT  3.805 1.795 4.035 2.125 ;
      RECT  3.805 2.125 8.515 2.355 ;
      RECT  4.925 2.355 5.155 2.675 ;
      RECT  6.045 2.355 6.275 2.675 ;
      RECT  7.165 2.355 7.395 2.675 ;
      RECT  8.285 2.355 8.515 2.675 ;
      RECT  3.805 2.355 4.035 3.245 ;
      RECT  3.805 3.245 4.3 3.475 ;
      RECT  1.72 4.365 2.76 4.595 ;
  END
END MDN_OR4B_4
#-----------------------------------------------------------------------
#      Cell        : MDN_TIE0_1
#      Description : Tie low
#      Equation    : X=0
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_TIE0_1
  CLASS CORE TIELOW ;
  FOREIGN MDN_TIE0_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.905 1.235 5.46 ;
      RECT  1.005 5.46 3.475 5.74 ;
      RECT  3.245 4.905 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.695 ;
      RECT  3.245 0.14 3.475 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 1.54 1.235 1.82 ;
    END
    ANTENNADIFFAREA 0.614 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.72 1.565 2.915 1.795 ;
      RECT  2.685 1.795 2.915 2.69 ;
      RECT  0.445 2.35 0.675 3.245 ;
      RECT  0.18 3.245 2.76 3.475 ;
      RECT  1.565 2.35 1.795 3.245 ;
  END
END MDN_TIE0_1
#-----------------------------------------------------------------------
#      Cell        : MDN_TIE1_1
#      Description : Tie high
#      Equation    : X=1
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_TIE1_1
  CLASS CORE TIEHIGH ;
  FOREIGN MDN_TIE1_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.48 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 4.905 1.235 5.46 ;
      RECT  1.005 5.46 3.475 5.74 ;
      RECT  3.245 4.905 3.475 5.46 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 4.48 5.74 ;
      LAYER VIA12 ;
      RECT  1.27 5.47 1.53 5.73 ;
      RECT  1.83 5.47 2.09 5.73 ;
      RECT  2.39 5.47 2.65 5.73 ;
      RECT  2.95 5.47 3.21 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  1.005 -0.14 3.475 0.14 ;
      RECT  1.005 0.14 1.235 0.695 ;
      RECT  3.245 0.14 3.475 0.695 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 4.48 0.14 ;
      LAYER VIA12 ;
      RECT  1.27 -0.13 1.53 0.13 ;
      RECT  1.83 -0.13 2.09 0.13 ;
      RECT  2.39 -0.13 2.65 0.13 ;
      RECT  2.95 -0.13 3.21 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.18 3.78 1.235 4.06 ;
    END
    ANTENNADIFFAREA 0.898 ;
  END X
  OBS
      LAYER METAL1 ;
      RECT  1.565 1.565 2.76 1.795 ;
      RECT  1.565 1.795 1.795 2.125 ;
      RECT  0.445 2.125 1.795 2.355 ;
      RECT  0.445 2.355 0.675 2.69 ;
      RECT  1.565 2.355 1.795 2.69 ;
      RECT  2.685 2.35 2.915 3.245 ;
      RECT  1.72 3.245 2.915 3.475 ;
  END
END MDN_TIE1_1
#-----------------------------------------------------------------------
#      Cell        : MDN_TIEDIP_1
#      Description : Antenna diode p+/nwell
#      Equation    : X=tristate(enable=0,data=0)
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_TIEDIP_1
  CLASS CORE ANTENNACELL ;
  FOREIGN MDN_TIEDIP_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.24 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 5.46 0.56 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 2.24 5.74 ;
      LAYER VIA12 ;
      RECT  0.15 5.47 0.41 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  -0.17 -0.14 0.56 0.14 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 2.24 0.14 ;
      LAYER VIA12 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  PIN X
    DIRECTION INOUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.445 3.78 1.29 4.06 ;
    END
    ANTENNADIFFAREA 1.472 ;
  END X
END MDN_TIEDIP_1

END LIBRARY
