#----------------------------------------------------------------------------
# Description	: Cell LEF definitions for ts18ugfsdmp
#		  (TSMC 018um fsg -StdVt Metal Programable Library)
# Date		: $Date: 2006/06/08 03:58:23 $
# Copyright	: 1997-2006 by Virage Logic Corporation
# Revision	: Version $Revision: 1.18 $
#----------------------------------------------------------------------------

VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

# Placement site definition for this library.
SITE ts18_dmp
  CLASS core ;
  SIZE 2.24 BY 5.6 ;
END ts18_dmp


#-----------------------------------------------------------------------
#      Cell        : MDN_FSDPQ_4
#      Description : D-Flip Flop w/scan, pos-edge triggered, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDPQ_4
  CLASS CORE ;
  FOREIGN MDN_FSDPQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.4 1.565 21.395 1.795 ;
      RECT  21.165 1.795 21.395 3.245 ;
      RECT  17.4 3.245 21.395 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 12.435 5.74 ;
      RECT  12.205 5.0 12.435 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.925 -0.14 19.6 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.36 -0.14 4.035 0.14 ;
      RECT  3.805 0.14 4.035 0.89 ;
      RECT  3.805 0.89 4.3 1.12 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  6.1 0.6 6.33 0.83 ;
      RECT  6.1 0.83 9.635 1.005 ;
      RECT  6.1 1.005 12.435 1.06 ;
      RECT  9.405 1.06 12.435 1.235 ;
      RECT  12.205 1.235 12.435 1.75 ;
      RECT  12.205 1.75 13.96 1.98 ;
      RECT  12.205 1.98 12.435 3.16 ;
      RECT  11.38 3.16 12.435 3.39 ;
      RECT  12.205 3.39 12.435 3.62 ;
      RECT  12.205 3.62 14.115 3.805 ;
      RECT  12.205 3.805 15.5 3.85 ;
      RECT  13.885 3.85 15.5 4.035 ;
      RECT  7.11 0.37 9.71 0.6 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.82 0.6 13.05 0.83 ;
      RECT  12.82 0.83 15.985 1.06 ;
      RECT  15.755 1.06 15.985 1.565 ;
      RECT  15.755 1.565 16.355 1.795 ;
      RECT  16.125 1.795 16.355 2.125 ;
      RECT  16.125 2.125 20.835 2.355 ;
      RECT  17.245 2.355 17.475 2.645 ;
      RECT  20.605 2.355 20.835 2.655 ;
      RECT  19.485 2.355 19.715 2.66 ;
      RECT  18.365 2.355 18.595 2.665 ;
      RECT  16.125 2.355 16.355 3.245 ;
      RECT  15.86 3.245 16.355 3.475 ;
      RECT  14.39 0.37 16.41 0.6 ;
      RECT  4.745 1.005 5.715 1.01 ;
      RECT  4.74 1.01 5.715 1.015 ;
      RECT  4.735 1.015 5.715 1.02 ;
      RECT  4.73 1.02 5.715 1.025 ;
      RECT  4.725 1.025 5.715 1.03 ;
      RECT  4.72 1.03 5.715 1.035 ;
      RECT  4.715 1.035 5.715 1.04 ;
      RECT  4.71 1.04 5.715 1.045 ;
      RECT  4.705 1.045 5.715 1.05 ;
      RECT  4.7 1.05 5.715 1.055 ;
      RECT  4.695 1.055 5.715 1.06 ;
      RECT  4.69 1.06 5.715 1.065 ;
      RECT  4.685 1.065 5.715 1.07 ;
      RECT  4.68 1.07 5.715 1.075 ;
      RECT  4.675 1.075 5.715 1.08 ;
      RECT  4.67 1.08 5.715 1.085 ;
      RECT  4.665 1.085 5.715 1.09 ;
      RECT  4.66 1.09 5.715 1.095 ;
      RECT  4.655 1.095 5.715 1.1 ;
      RECT  4.65 1.1 5.715 1.105 ;
      RECT  4.645 1.105 5.715 1.11 ;
      RECT  4.64 1.11 5.715 1.115 ;
      RECT  4.635 1.115 5.715 1.12 ;
      RECT  4.63 1.12 5.715 1.125 ;
      RECT  4.625 1.125 5.715 1.13 ;
      RECT  4.62 1.13 5.715 1.135 ;
      RECT  4.615 1.135 5.715 1.14 ;
      RECT  4.61 1.14 5.715 1.145 ;
      RECT  4.605 1.145 5.715 1.15 ;
      RECT  4.6 1.15 5.715 1.155 ;
      RECT  4.595 1.155 5.715 1.16 ;
      RECT  4.59 1.16 5.715 1.165 ;
      RECT  4.585 1.165 5.715 1.17 ;
      RECT  4.58 1.17 5.715 1.175 ;
      RECT  4.575 1.175 5.715 1.18 ;
      RECT  4.57 1.18 5.715 1.185 ;
      RECT  4.565 1.185 5.715 1.19 ;
      RECT  4.56 1.19 5.715 1.195 ;
      RECT  4.555 1.195 5.715 1.2 ;
      RECT  4.55 1.2 5.715 1.205 ;
      RECT  4.545 1.205 5.715 1.21 ;
      RECT  4.54 1.21 5.715 1.215 ;
      RECT  4.535 1.215 5.715 1.22 ;
      RECT  4.53 1.22 5.715 1.225 ;
      RECT  4.525 1.225 5.715 1.23 ;
      RECT  4.52 1.23 5.715 1.235 ;
      RECT  4.515 1.235 4.84 1.24 ;
      RECT  5.485 1.235 5.715 1.75 ;
      RECT  4.51 1.24 4.835 1.245 ;
      RECT  4.505 1.245 4.83 1.25 ;
      RECT  4.5 1.25 4.825 1.255 ;
      RECT  4.495 1.255 4.82 1.26 ;
      RECT  4.49 1.26 4.815 1.265 ;
      RECT  4.485 1.265 4.81 1.27 ;
      RECT  4.48 1.27 4.805 1.275 ;
      RECT  4.475 1.275 4.8 1.28 ;
      RECT  4.47 1.28 4.795 1.285 ;
      RECT  4.465 1.285 4.79 1.29 ;
      RECT  4.46 1.29 4.785 1.295 ;
      RECT  4.455 1.295 4.78 1.3 ;
      RECT  4.45 1.3 4.775 1.305 ;
      RECT  4.445 1.305 4.77 1.31 ;
      RECT  4.44 1.31 4.765 1.315 ;
      RECT  4.435 1.315 4.76 1.32 ;
      RECT  4.43 1.32 4.755 1.325 ;
      RECT  4.425 1.325 4.75 1.33 ;
      RECT  4.42 1.33 4.745 1.335 ;
      RECT  4.415 1.335 4.74 1.34 ;
      RECT  4.41 1.34 4.735 1.345 ;
      RECT  4.405 1.345 4.73 1.35 ;
      RECT  4.4 1.35 4.725 1.355 ;
      RECT  4.395 1.355 4.72 1.36 ;
      RECT  4.39 1.36 4.715 1.365 ;
      RECT  4.385 1.365 4.71 1.37 ;
      RECT  4.38 1.37 4.705 1.375 ;
      RECT  4.375 1.375 4.7 1.38 ;
      RECT  4.37 1.38 4.695 1.385 ;
      RECT  4.365 1.385 4.69 1.39 ;
      RECT  4.36 1.39 4.685 1.395 ;
      RECT  4.355 1.395 4.68 1.4 ;
      RECT  4.35 1.4 4.675 1.405 ;
      RECT  4.345 1.405 4.67 1.41 ;
      RECT  4.34 1.41 4.665 1.415 ;
      RECT  4.335 1.415 4.66 1.42 ;
      RECT  4.33 1.42 4.655 1.425 ;
      RECT  4.325 1.425 4.65 1.43 ;
      RECT  4.32 1.43 4.645 1.435 ;
      RECT  4.315 1.435 4.64 1.44 ;
      RECT  4.31 1.44 4.635 1.445 ;
      RECT  4.305 1.445 4.63 1.45 ;
      RECT  4.3 1.45 4.625 1.455 ;
      RECT  4.295 1.455 4.62 1.46 ;
      RECT  4.29 1.46 4.615 1.465 ;
      RECT  4.285 1.465 4.61 1.47 ;
      RECT  4.28 1.47 4.605 1.475 ;
      RECT  4.275 1.475 4.6 1.48 ;
      RECT  4.27 1.48 4.595 1.485 ;
      RECT  4.265 1.485 4.59 1.49 ;
      RECT  4.26 1.49 4.585 1.495 ;
      RECT  4.255 1.495 4.58 1.5 ;
      RECT  4.25 1.5 4.575 1.505 ;
      RECT  4.245 1.505 4.57 1.51 ;
      RECT  4.24 1.51 4.565 1.515 ;
      RECT  4.235 1.515 4.56 1.52 ;
      RECT  4.23 1.52 4.555 1.525 ;
      RECT  4.225 1.525 4.55 1.53 ;
      RECT  4.22 1.53 4.545 1.535 ;
      RECT  4.215 1.535 4.54 1.54 ;
      RECT  4.21 1.54 4.535 1.545 ;
      RECT  4.205 1.545 4.53 1.55 ;
      RECT  4.2 1.55 4.525 1.555 ;
      RECT  4.195 1.555 4.52 1.56 ;
      RECT  4.19 1.56 4.515 1.565 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  3.245 1.565 4.51 1.57 ;
      RECT  3.245 1.57 4.505 1.575 ;
      RECT  3.245 1.575 4.5 1.58 ;
      RECT  3.245 1.58 4.495 1.585 ;
      RECT  3.245 1.585 4.49 1.59 ;
      RECT  3.245 1.59 4.485 1.595 ;
      RECT  3.245 1.595 4.48 1.6 ;
      RECT  3.245 1.6 4.475 1.605 ;
      RECT  3.245 1.605 4.47 1.61 ;
      RECT  3.245 1.61 4.465 1.615 ;
      RECT  3.245 1.615 4.46 1.62 ;
      RECT  3.245 1.62 4.455 1.625 ;
      RECT  3.245 1.625 4.45 1.63 ;
      RECT  3.245 1.63 4.445 1.635 ;
      RECT  3.245 1.635 4.44 1.64 ;
      RECT  3.245 1.64 4.435 1.645 ;
      RECT  3.245 1.645 4.43 1.65 ;
      RECT  3.245 1.65 4.425 1.655 ;
      RECT  3.245 1.655 4.42 1.66 ;
      RECT  3.245 1.66 4.415 1.665 ;
      RECT  3.245 1.665 4.41 1.67 ;
      RECT  3.245 1.67 4.405 1.675 ;
      RECT  3.245 1.675 4.4 1.68 ;
      RECT  3.245 1.68 4.395 1.685 ;
      RECT  3.245 1.685 4.39 1.69 ;
      RECT  3.245 1.69 4.385 1.695 ;
      RECT  3.245 1.695 4.38 1.7 ;
      RECT  3.245 1.7 4.375 1.705 ;
      RECT  3.245 1.705 4.37 1.71 ;
      RECT  3.245 1.71 4.365 1.715 ;
      RECT  3.245 1.715 4.36 1.72 ;
      RECT  3.245 1.72 4.355 1.725 ;
      RECT  3.245 1.725 4.35 1.73 ;
      RECT  3.245 1.73 4.345 1.735 ;
      RECT  3.245 1.735 4.34 1.74 ;
      RECT  3.245 1.74 4.335 1.745 ;
      RECT  3.245 1.745 4.33 1.75 ;
      RECT  3.245 1.75 4.325 1.755 ;
      RECT  5.485 1.75 7.24 1.98 ;
      RECT  3.245 1.755 4.32 1.76 ;
      RECT  3.245 1.76 4.315 1.765 ;
      RECT  3.245 1.765 4.31 1.77 ;
      RECT  3.245 1.77 4.305 1.775 ;
      RECT  3.245 1.775 4.3 1.78 ;
      RECT  3.245 1.78 4.295 1.785 ;
      RECT  3.245 1.785 4.29 1.79 ;
      RECT  3.245 1.79 4.285 1.795 ;
      RECT  6.2 1.29 8.78 1.52 ;
      RECT  12.92 1.29 15.5 1.52 ;
      RECT  9.965 1.565 11.02 1.795 ;
      RECT  9.965 1.795 10.195 2.405 ;
      RECT  9.35 2.405 10.195 2.635 ;
      RECT  9.965 2.635 10.195 3.755 ;
      RECT  9.965 3.755 11.875 3.985 ;
      RECT  11.645 3.985 11.875 4.08 ;
      RECT  11.645 4.08 13.555 4.31 ;
      RECT  13.325 4.31 13.555 4.365 ;
      RECT  13.325 4.365 14.675 4.595 ;
      RECT  14.445 4.595 14.675 4.995 ;
      RECT  14.445 4.995 15.19 5.0 ;
      RECT  14.445 5.0 15.29 5.225 ;
      RECT  14.95 5.225 15.29 5.23 ;
      RECT  4.66 1.75 5.155 1.98 ;
      RECT  4.925 1.98 5.155 2.405 ;
      RECT  3.75 2.405 5.155 2.635 ;
      RECT  4.925 2.635 5.155 3.245 ;
      RECT  4.66 3.245 5.155 3.475 ;
      RECT  7.67 1.75 8.01 1.98 ;
      RECT  7.725 1.98 7.955 3.435 ;
      RECT  8.285 1.75 9.48 1.98 ;
      RECT  8.285 1.98 8.515 3.245 ;
      RECT  8.285 3.245 9.37 3.475 ;
      RECT  9.14 3.475 9.37 4.215 ;
      RECT  9.14 4.215 11.315 4.445 ;
      RECT  11.085 4.445 11.315 4.54 ;
      RECT  11.085 4.54 12.995 4.77 ;
      RECT  12.765 4.77 12.995 5.0 ;
      RECT  12.765 5.0 14.17 5.23 ;
      RECT  14.39 1.75 14.73 1.98 ;
      RECT  14.445 1.98 14.675 3.53 ;
      RECT  12.92 3.16 13.98 3.39 ;
      RECT  6.2 3.245 7.24 3.475 ;
      RECT  1.72 3.805 2.76 4.035 ;
      RECT  3.19 3.805 8.78 4.035 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  9.405 4.675 10.755 4.905 ;
      RECT  9.405 4.905 9.635 4.925 ;
      RECT  10.525 4.905 10.755 5.0 ;
      RECT  7.67 4.925 9.635 5.155 ;
      RECT  10.525 5.0 11.93 5.23 ;
      RECT  1.51 5.0 5.21 5.23 ;
  END
END MDN_FSDPQ_4
