#----------------------------------------------------------------------------
# Description	: Cell LEF definitions for ts18ugfsdmp
#		  (TSMC 018um fsg -StdVt Metal Programable Library)
# Date		: $Date: 2006/06/08 03:58:23 $
# Copyright	: 1997-2006 by Virage Logic Corporation
# Revision	: Version $Revision: 1.18 $
#----------------------------------------------------------------------------

VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

# Placement site definition for this library.
SITE ts18_dmp
  CLASS core ;
  SIZE 2.24 BY 5.6 ;
END ts18_dmp



#-----------------------------------------------------------------------
#      Cell        : MDN_FSDPQ_4
#      Description : D-Flip Flop w/scan, pos-edge triggered, q-only
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDPQ_4
  CLASS CORE ;
  FOREIGN MDN_FSDPQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.4 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  10.5 2.125 10.78 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 2.125 2.94 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  17.4 1.565 21.395 1.795 ;
      RECT  21.165 1.795 21.395 3.245 ;
      RECT  17.4 3.245 21.395 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  21.165 5.46 22.57 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.925 5.46 19.6 5.74 ;
      RECT  16.685 4.9 16.915 5.46 ;
      RECT  16.685 5.46 17.36 5.74 ;
      RECT  9.91 5.135 10.25 5.46 ;
      RECT  9.52 5.46 12.435 5.74 ;
      RECT  12.205 5.0 12.435 5.46 ;
      RECT  5.485 4.9 5.715 5.46 ;
      RECT  5.04 5.46 5.715 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 22.4 5.74 ;
      LAYER VIA12 ;
      RECT  21.43 5.47 21.69 5.73 ;
      RECT  21.99 5.47 22.25 5.73 ;
      RECT  19.19 5.47 19.45 5.73 ;
      RECT  16.95 5.47 17.21 5.73 ;
      RECT  9.67 5.47 9.93 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  10.79 5.47 11.05 5.73 ;
      RECT  11.35 5.47 11.61 5.73 ;
      RECT  11.91 5.47 12.17 5.73 ;
      RECT  5.19 5.47 5.45 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  21.165 -0.14 22.57 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  18.925 -0.14 19.6 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  16.24 -0.14 16.915 0.14 ;
      RECT  16.685 0.14 16.915 0.7 ;
      RECT  9.965 -0.14 12.435 0.14 ;
      RECT  9.965 0.14 10.195 0.73 ;
      RECT  12.205 0.14 12.435 0.73 ;
      RECT  5.485 -0.14 6.16 0.14 ;
      RECT  5.485 0.14 5.715 0.73 ;
      RECT  3.36 -0.14 4.035 0.14 ;
      RECT  3.805 0.14 4.035 0.89 ;
      RECT  3.805 0.89 4.3 1.12 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 22.4 0.14 ;
      LAYER VIA12 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  16.39 -0.13 16.65 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  11.35 -0.13 11.61 0.13 ;
      RECT  11.91 -0.13 12.17 0.13 ;
      RECT  5.75 -0.13 6.01 0.13 ;
      RECT  3.51 -0.13 3.77 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.99 0.37 6.33 0.6 ;
      RECT  6.1 0.6 6.33 0.83 ;
      RECT  6.1 0.83 9.635 1.005 ;
      RECT  6.1 1.005 12.435 1.06 ;
      RECT  9.405 1.06 12.435 1.235 ;
      RECT  12.205 1.235 12.435 1.75 ;
      RECT  12.205 1.75 13.96 1.98 ;
      RECT  12.205 1.98 12.435 3.16 ;
      RECT  11.38 3.16 12.435 3.39 ;
      RECT  12.205 3.39 12.435 3.62 ;
      RECT  12.205 3.62 14.115 3.805 ;
      RECT  12.205 3.805 15.5 3.85 ;
      RECT  13.885 3.85 15.5 4.035 ;
      RECT  7.11 0.37 9.71 0.6 ;
      RECT  12.71 0.37 13.05 0.6 ;
      RECT  12.82 0.6 13.05 0.83 ;
      RECT  12.82 0.83 15.985 1.06 ;
      RECT  15.755 1.06 15.985 1.565 ;
      RECT  15.755 1.565 16.355 1.795 ;
      RECT  16.125 1.795 16.355 2.125 ;
      RECT  16.125 2.125 20.835 2.355 ;
      RECT  17.245 2.355 17.475 2.645 ;
      RECT  20.605 2.355 20.835 2.655 ;
      RECT  19.485 2.355 19.715 2.66 ;
      RECT  18.365 2.355 18.595 2.665 ;
      RECT  16.125 2.355 16.355 3.245 ;
      RECT  15.86 3.245 16.355 3.475 ;
      RECT  14.39 0.37 16.41 0.6 ;
      RECT  4.745 1.005 5.715 1.01 ;
      RECT  4.74 1.01 5.715 1.015 ;
      RECT  4.735 1.015 5.715 1.02 ;
      RECT  4.73 1.02 5.715 1.025 ;
      RECT  4.725 1.025 5.715 1.03 ;
      RECT  4.72 1.03 5.715 1.035 ;
      RECT  4.715 1.035 5.715 1.04 ;
      RECT  4.71 1.04 5.715 1.045 ;
      RECT  4.705 1.045 5.715 1.05 ;
      RECT  4.7 1.05 5.715 1.055 ;
      RECT  4.695 1.055 5.715 1.06 ;
      RECT  4.69 1.06 5.715 1.065 ;
      RECT  4.685 1.065 5.715 1.07 ;
      RECT  4.68 1.07 5.715 1.075 ;
      RECT  4.675 1.075 5.715 1.08 ;
      RECT  4.67 1.08 5.715 1.085 ;
      RECT  4.665 1.085 5.715 1.09 ;
      RECT  4.66 1.09 5.715 1.095 ;
      RECT  4.655 1.095 5.715 1.1 ;
      RECT  4.65 1.1 5.715 1.105 ;
      RECT  4.645 1.105 5.715 1.11 ;
      RECT  4.64 1.11 5.715 1.115 ;
      RECT  4.635 1.115 5.715 1.12 ;
      RECT  4.63 1.12 5.715 1.125 ;
      RECT  4.625 1.125 5.715 1.13 ;
      RECT  4.62 1.13 5.715 1.135 ;
      RECT  4.615 1.135 5.715 1.14 ;
      RECT  4.61 1.14 5.715 1.145 ;
      RECT  4.605 1.145 5.715 1.15 ;
      RECT  4.6 1.15 5.715 1.155 ;
      RECT  4.595 1.155 5.715 1.16 ;
      RECT  4.59 1.16 5.715 1.165 ;
      RECT  4.585 1.165 5.715 1.17 ;
      RECT  4.58 1.17 5.715 1.175 ;
      RECT  4.575 1.175 5.715 1.18 ;
      RECT  4.57 1.18 5.715 1.185 ;
      RECT  4.565 1.185 5.715 1.19 ;
      RECT  4.56 1.19 5.715 1.195 ;
      RECT  4.555 1.195 5.715 1.2 ;
      RECT  4.55 1.2 5.715 1.205 ;
      RECT  4.545 1.205 5.715 1.21 ;
      RECT  4.54 1.21 5.715 1.215 ;
      RECT  4.535 1.215 5.715 1.22 ;
      RECT  4.53 1.22 5.715 1.225 ;
      RECT  4.525 1.225 5.715 1.23 ;
      RECT  4.52 1.23 5.715 1.235 ;
      RECT  4.515 1.235 4.84 1.24 ;
      RECT  5.485 1.235 5.715 1.75 ;
      RECT  4.51 1.24 4.835 1.245 ;
      RECT  4.505 1.245 4.83 1.25 ;
      RECT  4.5 1.25 4.825 1.255 ;
      RECT  4.495 1.255 4.82 1.26 ;
      RECT  4.49 1.26 4.815 1.265 ;
      RECT  4.485 1.265 4.81 1.27 ;
      RECT  4.48 1.27 4.805 1.275 ;
      RECT  4.475 1.275 4.8 1.28 ;
      RECT  4.47 1.28 4.795 1.285 ;
      RECT  4.465 1.285 4.79 1.29 ;
      RECT  4.46 1.29 4.785 1.295 ;
      RECT  4.455 1.295 4.78 1.3 ;
      RECT  4.45 1.3 4.775 1.305 ;
      RECT  4.445 1.305 4.77 1.31 ;
      RECT  4.44 1.31 4.765 1.315 ;
      RECT  4.435 1.315 4.76 1.32 ;
      RECT  4.43 1.32 4.755 1.325 ;
      RECT  4.425 1.325 4.75 1.33 ;
      RECT  4.42 1.33 4.745 1.335 ;
      RECT  4.415 1.335 4.74 1.34 ;
      RECT  4.41 1.34 4.735 1.345 ;
      RECT  4.405 1.345 4.73 1.35 ;
      RECT  4.4 1.35 4.725 1.355 ;
      RECT  4.395 1.355 4.72 1.36 ;
      RECT  4.39 1.36 4.715 1.365 ;
      RECT  4.385 1.365 4.71 1.37 ;
      RECT  4.38 1.37 4.705 1.375 ;
      RECT  4.375 1.375 4.7 1.38 ;
      RECT  4.37 1.38 4.695 1.385 ;
      RECT  4.365 1.385 4.69 1.39 ;
      RECT  4.36 1.39 4.685 1.395 ;
      RECT  4.355 1.395 4.68 1.4 ;
      RECT  4.35 1.4 4.675 1.405 ;
      RECT  4.345 1.405 4.67 1.41 ;
      RECT  4.34 1.41 4.665 1.415 ;
      RECT  4.335 1.415 4.66 1.42 ;
      RECT  4.33 1.42 4.655 1.425 ;
      RECT  4.325 1.425 4.65 1.43 ;
      RECT  4.32 1.43 4.645 1.435 ;
      RECT  4.315 1.435 4.64 1.44 ;
      RECT  4.31 1.44 4.635 1.445 ;
      RECT  4.305 1.445 4.63 1.45 ;
      RECT  4.3 1.45 4.625 1.455 ;
      RECT  4.295 1.455 4.62 1.46 ;
      RECT  4.29 1.46 4.615 1.465 ;
      RECT  4.285 1.465 4.61 1.47 ;
      RECT  4.28 1.47 4.605 1.475 ;
      RECT  4.275 1.475 4.6 1.48 ;
      RECT  4.27 1.48 4.595 1.485 ;
      RECT  4.265 1.485 4.59 1.49 ;
      RECT  4.26 1.49 4.585 1.495 ;
      RECT  4.255 1.495 4.58 1.5 ;
      RECT  4.25 1.5 4.575 1.505 ;
      RECT  4.245 1.505 4.57 1.51 ;
      RECT  4.24 1.51 4.565 1.515 ;
      RECT  4.235 1.515 4.56 1.52 ;
      RECT  4.23 1.52 4.555 1.525 ;
      RECT  4.225 1.525 4.55 1.53 ;
      RECT  4.22 1.53 4.545 1.535 ;
      RECT  4.215 1.535 4.54 1.54 ;
      RECT  4.21 1.54 4.535 1.545 ;
      RECT  4.205 1.545 4.53 1.55 ;
      RECT  4.2 1.55 4.525 1.555 ;
      RECT  4.195 1.555 4.52 1.56 ;
      RECT  4.19 1.56 4.515 1.565 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  3.245 1.565 4.51 1.57 ;
      RECT  3.245 1.57 4.505 1.575 ;
      RECT  3.245 1.575 4.5 1.58 ;
      RECT  3.245 1.58 4.495 1.585 ;
      RECT  3.245 1.585 4.49 1.59 ;
      RECT  3.245 1.59 4.485 1.595 ;
      RECT  3.245 1.595 4.48 1.6 ;
      RECT  3.245 1.6 4.475 1.605 ;
      RECT  3.245 1.605 4.47 1.61 ;
      RECT  3.245 1.61 4.465 1.615 ;
      RECT  3.245 1.615 4.46 1.62 ;
      RECT  3.245 1.62 4.455 1.625 ;
      RECT  3.245 1.625 4.45 1.63 ;
      RECT  3.245 1.63 4.445 1.635 ;
      RECT  3.245 1.635 4.44 1.64 ;
      RECT  3.245 1.64 4.435 1.645 ;
      RECT  3.245 1.645 4.43 1.65 ;
      RECT  3.245 1.65 4.425 1.655 ;
      RECT  3.245 1.655 4.42 1.66 ;
      RECT  3.245 1.66 4.415 1.665 ;
      RECT  3.245 1.665 4.41 1.67 ;
      RECT  3.245 1.67 4.405 1.675 ;
      RECT  3.245 1.675 4.4 1.68 ;
      RECT  3.245 1.68 4.395 1.685 ;
      RECT  3.245 1.685 4.39 1.69 ;
      RECT  3.245 1.69 4.385 1.695 ;
      RECT  3.245 1.695 4.38 1.7 ;
      RECT  3.245 1.7 4.375 1.705 ;
      RECT  3.245 1.705 4.37 1.71 ;
      RECT  3.245 1.71 4.365 1.715 ;
      RECT  3.245 1.715 4.36 1.72 ;
      RECT  3.245 1.72 4.355 1.725 ;
      RECT  3.245 1.725 4.35 1.73 ;
      RECT  3.245 1.73 4.345 1.735 ;
      RECT  3.245 1.735 4.34 1.74 ;
      RECT  3.245 1.74 4.335 1.745 ;
      RECT  3.245 1.745 4.33 1.75 ;
      RECT  3.245 1.75 4.325 1.755 ;
      RECT  5.485 1.75 7.24 1.98 ;
      RECT  3.245 1.755 4.32 1.76 ;
      RECT  3.245 1.76 4.315 1.765 ;
      RECT  3.245 1.765 4.31 1.77 ;
      RECT  3.245 1.77 4.305 1.775 ;
      RECT  3.245 1.775 4.3 1.78 ;
      RECT  3.245 1.78 4.295 1.785 ;
      RECT  3.245 1.785 4.29 1.79 ;
      RECT  3.245 1.79 4.285 1.795 ;
      RECT  6.2 1.29 8.78 1.52 ;
      RECT  12.92 1.29 15.5 1.52 ;
      RECT  9.965 1.565 11.02 1.795 ;
      RECT  9.965 1.795 10.195 2.405 ;
      RECT  9.35 2.405 10.195 2.635 ;
      RECT  9.965 2.635 10.195 3.755 ;
      RECT  9.965 3.755 11.875 3.985 ;
      RECT  11.645 3.985 11.875 4.08 ;
      RECT  11.645 4.08 13.555 4.31 ;
      RECT  13.325 4.31 13.555 4.365 ;
      RECT  13.325 4.365 14.675 4.595 ;
      RECT  14.445 4.595 14.675 4.995 ;
      RECT  14.445 4.995 15.19 5.0 ;
      RECT  14.445 5.0 15.29 5.225 ;
      RECT  14.95 5.225 15.29 5.23 ;
      RECT  4.66 1.75 5.155 1.98 ;
      RECT  4.925 1.98 5.155 2.405 ;
      RECT  3.75 2.405 5.155 2.635 ;
      RECT  4.925 2.635 5.155 3.245 ;
      RECT  4.66 3.245 5.155 3.475 ;
      RECT  7.67 1.75 8.01 1.98 ;
      RECT  7.725 1.98 7.955 3.435 ;
      RECT  8.285 1.75 9.48 1.98 ;
      RECT  8.285 1.98 8.515 3.245 ;
      RECT  8.285 3.245 9.37 3.475 ;
      RECT  9.14 3.475 9.37 4.215 ;
      RECT  9.14 4.215 11.315 4.445 ;
      RECT  11.085 4.445 11.315 4.54 ;
      RECT  11.085 4.54 12.995 4.77 ;
      RECT  12.765 4.77 12.995 5.0 ;
      RECT  12.765 5.0 14.17 5.23 ;
      RECT  14.39 1.75 14.73 1.98 ;
      RECT  14.445 1.98 14.675 3.53 ;
      RECT  12.92 3.16 13.98 3.39 ;
      RECT  6.2 3.245 7.24 3.475 ;
      RECT  1.72 3.805 2.76 4.035 ;
      RECT  3.19 3.805 8.78 4.035 ;
      RECT  0.18 4.365 4.3 4.595 ;
      RECT  9.405 4.675 10.755 4.905 ;
      RECT  9.405 4.905 9.635 4.925 ;
      RECT  10.525 4.905 10.755 5.0 ;
      RECT  7.67 4.925 9.635 5.155 ;
      RECT  10.525 5.0 11.93 5.23 ;
      RECT  1.51 5.0 5.21 5.23 ;
  END
END MDN_FSDPQ_4

#-----------------------------------------------------------------------
#      Cell        : MDN_FSDPRB_4
#      Description : D-Flip Flop w/scan, pos-edge triggered, lo-async-clear
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq:QN=iqn
#      Version     : $Revision: 1.18 $
#      Created     : $Date: 2006/06/08 03:58:23 $
#
MACRO MDN_FSDPRB_4
  CLASS CORE ;
  FOREIGN MDN_FSDPRB_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 29.12 BY 5.6 ;
  SYMMETRY  X ;
  SITE ts18_dmp ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  4.9 2.125 5.18 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  2.66 1.565 2.94 2.69 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  19.64 1.565 22.92 1.795 ;
      RECT  22.285 1.795 22.515 3.245 ;
      RECT  19.64 3.245 22.92 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER METAL1 ;
      RECT  24.82 1.565 28.94 1.795 ;
      RECT  26.765 1.795 26.995 3.245 ;
      RECT  24.82 3.245 28.94 3.475 ;
    END
    ANTENNADIFFAREA 6.048 ;
  END QN
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  14.98 2.125 16.38 2.355 ;
      RECT  14.98 2.355 15.26 2.915 ;
      RECT  16.1 2.355 16.38 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  1.54 2.125 1.82 2.915 ;
    END
    ANTENNAGATEAREA 1.134 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER METAL1 ;
      RECT  0.42 2.125 0.7 2.915 ;
    END
    ANTENNAGATEAREA 0.567 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  27.885 4.9 28.115 5.46 ;
      RECT  27.885 5.46 29.29 5.74 ;
      RECT  25.645 4.9 25.875 5.46 ;
      RECT  25.645 5.46 26.32 5.74 ;
      RECT  23.405 4.9 23.635 5.46 ;
      RECT  23.405 5.46 24.08 5.74 ;
      RECT  21.165 4.9 21.395 5.46 ;
      RECT  20.72 5.46 21.395 5.74 ;
      RECT  18.925 4.9 19.155 5.46 ;
      RECT  18.48 5.46 19.155 5.74 ;
      RECT  14.445 5.08 14.675 5.46 ;
      RECT  14.445 5.46 16.915 5.74 ;
      RECT  16.685 4.93 16.915 5.46 ;
      RECT  9.965 5.08 10.195 5.46 ;
      RECT  9.965 5.46 10.64 5.74 ;
      RECT  5.485 5.0 5.715 5.46 ;
      RECT  5.485 5.46 6.16 5.74 ;
      RECT  1.005 4.87 1.235 5.46 ;
      RECT  -0.17 5.46 1.235 5.74 ;
      LAYER METAL2 ;
      RECT  0.0 5.46 29.12 5.74 ;
      LAYER VIA12 ;
      RECT  28.15 5.47 28.41 5.73 ;
      RECT  28.71 5.47 28.97 5.73 ;
      RECT  25.91 5.47 26.17 5.73 ;
      RECT  23.67 5.47 23.93 5.73 ;
      RECT  20.87 5.47 21.13 5.73 ;
      RECT  18.63 5.47 18.89 5.73 ;
      RECT  14.71 5.47 14.97 5.73 ;
      RECT  15.27 5.47 15.53 5.73 ;
      RECT  15.83 5.47 16.09 5.73 ;
      RECT  16.39 5.47 16.65 5.73 ;
      RECT  10.23 5.47 10.49 5.73 ;
      RECT  5.75 5.47 6.01 5.73 ;
      RECT  0.15 5.47 0.41 5.73 ;
      RECT  0.71 5.47 0.97 5.73 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
      RECT  25.645 -0.14 29.29 0.14 ;
      RECT  25.645 0.14 25.875 0.7 ;
      RECT  27.885 0.14 28.115 0.7 ;
      RECT  21.165 -0.14 23.635 0.14 ;
      RECT  21.165 0.14 21.395 0.7 ;
      RECT  23.405 0.14 23.635 0.73 ;
      RECT  18.925 -0.14 19.6 0.14 ;
      RECT  18.925 0.14 19.155 0.7 ;
      RECT  15.12 -0.14 16.24 0.14 ;
      RECT  15.565 0.14 15.795 0.89 ;
      RECT  15.16 0.89 16.2 1.12 ;
      RECT  9.965 -0.14 11.37 0.14 ;
      RECT  9.965 0.14 10.195 0.6 ;
      RECT  3.805 -0.14 5.715 0.14 ;
      RECT  5.485 0.14 5.715 0.6 ;
      RECT  3.805 0.14 4.035 1.005 ;
      RECT  3.805 1.005 4.3 1.235 ;
      RECT  -0.17 -0.14 0.675 0.14 ;
      RECT  0.445 0.14 0.675 1.005 ;
      RECT  0.18 1.005 0.675 1.235 ;
      LAYER METAL2 ;
      RECT  0.0 -0.14 29.12 0.14 ;
      LAYER VIA12 ;
      RECT  25.91 -0.13 26.17 0.13 ;
      RECT  26.47 -0.13 26.73 0.13 ;
      RECT  27.03 -0.13 27.29 0.13 ;
      RECT  27.59 -0.13 27.85 0.13 ;
      RECT  28.15 -0.13 28.41 0.13 ;
      RECT  28.71 -0.13 28.97 0.13 ;
      RECT  21.43 -0.13 21.69 0.13 ;
      RECT  21.99 -0.13 22.25 0.13 ;
      RECT  22.55 -0.13 22.81 0.13 ;
      RECT  23.11 -0.13 23.37 0.13 ;
      RECT  19.19 -0.13 19.45 0.13 ;
      RECT  15.27 -0.13 15.53 0.13 ;
      RECT  15.83 -0.13 16.09 0.13 ;
      RECT  10.23 -0.13 10.49 0.13 ;
      RECT  10.79 -0.13 11.05 0.13 ;
      RECT  4.07 -0.13 4.33 0.13 ;
      RECT  4.63 -0.13 4.89 0.13 ;
      RECT  5.19 -0.13 5.45 0.13 ;
      RECT  0.15 -0.13 0.41 0.13 ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
      RECT  5.98 0.37 6.33 0.6 ;
      RECT  5.98 0.6 6.21 0.83 ;
      RECT  4.715 0.83 6.21 1.06 ;
      RECT  4.715 1.06 4.945 1.29 ;
      RECT  10.425 0.37 13.05 0.6 ;
      RECT  10.425 0.6 10.655 0.83 ;
      RECT  7.11 0.37 9.635 0.6 ;
      RECT  9.405 0.6 9.635 0.83 ;
      RECT  9.405 0.83 10.655 1.06 ;
      RECT  23.91 0.37 24.25 0.6 ;
      RECT  23.91 0.6 24.14 1.005 ;
      RECT  21.67 0.37 23.13 0.6 ;
      RECT  22.9 0.6 23.13 1.005 ;
      RECT  22.9 1.005 24.14 1.235 ;
      RECT  26.15 0.37 27.61 0.6 ;
      RECT  6.44 0.83 8.78 1.06 ;
      RECT  8.44 1.06 8.78 1.12 ;
      RECT  6.44 1.06 6.67 1.29 ;
      RECT  5.485 1.29 6.67 1.52 ;
      RECT  5.485 1.52 5.715 1.565 ;
      RECT  1.72 1.005 3.475 1.235 ;
      RECT  3.245 1.235 3.475 1.565 ;
      RECT  3.245 1.565 5.715 1.795 ;
      RECT  10.905 0.83 13.96 1.06 ;
      RECT  13.62 1.06 13.96 1.12 ;
      RECT  10.905 1.06 11.135 1.29 ;
      RECT  8.94 1.29 11.135 1.295 ;
      RECT  8.935 1.295 11.135 1.3 ;
      RECT  8.93 1.3 11.135 1.305 ;
      RECT  8.925 1.305 11.135 1.31 ;
      RECT  8.92 1.31 11.135 1.315 ;
      RECT  8.915 1.315 11.135 1.32 ;
      RECT  8.91 1.32 11.135 1.325 ;
      RECT  8.905 1.325 11.135 1.33 ;
      RECT  8.9 1.33 11.135 1.335 ;
      RECT  8.895 1.335 11.135 1.34 ;
      RECT  8.89 1.34 11.135 1.345 ;
      RECT  8.885 1.345 11.135 1.35 ;
      RECT  8.88 1.35 11.135 1.355 ;
      RECT  8.875 1.355 11.135 1.36 ;
      RECT  8.87 1.36 11.135 1.365 ;
      RECT  8.865 1.365 11.135 1.37 ;
      RECT  8.86 1.37 11.135 1.375 ;
      RECT  8.855 1.375 11.135 1.38 ;
      RECT  8.85 1.38 11.135 1.385 ;
      RECT  8.845 1.385 11.135 1.39 ;
      RECT  8.84 1.39 11.135 1.395 ;
      RECT  8.835 1.395 11.135 1.4 ;
      RECT  8.83 1.4 11.135 1.405 ;
      RECT  8.825 1.405 11.135 1.41 ;
      RECT  8.82 1.41 11.135 1.415 ;
      RECT  8.815 1.415 11.135 1.42 ;
      RECT  6.9 1.29 8.215 1.295 ;
      RECT  6.9 1.295 8.22 1.3 ;
      RECT  6.9 1.3 8.225 1.305 ;
      RECT  6.9 1.305 8.23 1.31 ;
      RECT  6.9 1.31 8.235 1.315 ;
      RECT  6.9 1.315 8.24 1.32 ;
      RECT  6.9 1.32 8.245 1.325 ;
      RECT  6.9 1.325 8.25 1.33 ;
      RECT  6.9 1.33 8.255 1.335 ;
      RECT  6.9 1.335 8.26 1.34 ;
      RECT  6.9 1.34 8.265 1.345 ;
      RECT  6.9 1.345 8.27 1.35 ;
      RECT  6.9 1.35 8.275 1.355 ;
      RECT  6.9 1.355 8.28 1.36 ;
      RECT  6.9 1.36 8.285 1.365 ;
      RECT  6.9 1.365 8.29 1.37 ;
      RECT  6.9 1.37 8.295 1.375 ;
      RECT  6.9 1.375 8.3 1.38 ;
      RECT  6.9 1.38 8.305 1.385 ;
      RECT  6.9 1.385 8.31 1.39 ;
      RECT  6.9 1.39 8.315 1.395 ;
      RECT  6.9 1.395 8.32 1.4 ;
      RECT  6.9 1.4 8.325 1.405 ;
      RECT  6.9 1.405 8.33 1.41 ;
      RECT  6.9 1.41 8.335 1.415 ;
      RECT  6.9 1.415 8.34 1.42 ;
      RECT  6.9 1.42 11.135 1.52 ;
      RECT  8.11 1.52 9.035 1.525 ;
      RECT  8.115 1.525 9.03 1.53 ;
      RECT  8.12 1.53 9.025 1.535 ;
      RECT  8.125 1.535 9.02 1.54 ;
      RECT  8.13 1.54 9.015 1.545 ;
      RECT  8.135 1.545 9.01 1.55 ;
      RECT  8.14 1.55 9.005 1.555 ;
      RECT  8.145 1.555 9.0 1.56 ;
      RECT  8.15 1.56 8.995 1.565 ;
      RECT  8.155 1.565 8.99 1.57 ;
      RECT  8.16 1.57 8.985 1.575 ;
      RECT  8.165 1.575 8.98 1.58 ;
      RECT  8.17 1.58 8.975 1.585 ;
      RECT  8.175 1.585 8.97 1.59 ;
      RECT  8.18 1.59 8.965 1.595 ;
      RECT  8.185 1.595 8.96 1.6 ;
      RECT  8.19 1.6 8.955 1.605 ;
      RECT  8.195 1.605 8.95 1.61 ;
      RECT  8.2 1.61 8.945 1.615 ;
      RECT  8.205 1.615 8.94 1.62 ;
      RECT  8.21 1.62 8.935 1.625 ;
      RECT  8.215 1.625 8.93 1.63 ;
      RECT  8.22 1.63 8.925 1.635 ;
      RECT  8.225 1.635 8.92 1.64 ;
      RECT  8.23 1.64 8.915 1.645 ;
      RECT  8.235 1.645 8.91 1.65 ;
      RECT  16.685 1.005 18.445 1.235 ;
      RECT  16.685 1.235 16.915 1.565 ;
      RECT  11.38 1.29 13.465 1.295 ;
      RECT  11.38 1.295 13.47 1.3 ;
      RECT  11.38 1.3 13.475 1.305 ;
      RECT  11.38 1.305 13.48 1.31 ;
      RECT  11.38 1.31 13.485 1.315 ;
      RECT  11.38 1.315 13.49 1.32 ;
      RECT  11.38 1.32 13.495 1.325 ;
      RECT  11.38 1.325 13.5 1.33 ;
      RECT  11.38 1.33 13.505 1.335 ;
      RECT  11.38 1.335 13.51 1.34 ;
      RECT  11.38 1.34 13.515 1.345 ;
      RECT  11.38 1.345 13.52 1.35 ;
      RECT  11.38 1.35 13.525 1.355 ;
      RECT  11.38 1.355 13.53 1.36 ;
      RECT  11.38 1.36 13.535 1.365 ;
      RECT  11.38 1.365 13.54 1.37 ;
      RECT  11.38 1.37 13.545 1.375 ;
      RECT  11.38 1.375 13.55 1.38 ;
      RECT  11.38 1.38 13.555 1.385 ;
      RECT  11.38 1.385 13.56 1.39 ;
      RECT  11.38 1.39 13.565 1.395 ;
      RECT  11.38 1.395 13.57 1.4 ;
      RECT  11.38 1.4 13.575 1.405 ;
      RECT  11.38 1.405 13.58 1.41 ;
      RECT  11.38 1.41 13.585 1.415 ;
      RECT  11.38 1.415 13.59 1.42 ;
      RECT  11.38 1.42 13.595 1.425 ;
      RECT  11.38 1.425 13.6 1.43 ;
      RECT  11.38 1.43 13.605 1.435 ;
      RECT  11.38 1.435 13.61 1.44 ;
      RECT  11.38 1.44 13.615 1.445 ;
      RECT  11.38 1.445 13.62 1.45 ;
      RECT  11.38 1.45 13.625 1.455 ;
      RECT  11.38 1.455 13.63 1.46 ;
      RECT  11.38 1.46 13.635 1.465 ;
      RECT  11.38 1.465 13.64 1.47 ;
      RECT  11.38 1.47 13.645 1.475 ;
      RECT  11.38 1.475 13.65 1.48 ;
      RECT  11.38 1.48 13.655 1.485 ;
      RECT  11.38 1.485 13.66 1.49 ;
      RECT  11.38 1.49 13.665 1.495 ;
      RECT  11.38 1.495 13.67 1.5 ;
      RECT  11.38 1.5 13.675 1.505 ;
      RECT  11.38 1.505 13.68 1.51 ;
      RECT  11.38 1.51 13.685 1.515 ;
      RECT  11.38 1.515 13.69 1.52 ;
      RECT  13.36 1.52 13.695 1.525 ;
      RECT  13.365 1.525 13.7 1.53 ;
      RECT  13.37 1.53 13.705 1.535 ;
      RECT  13.375 1.535 13.71 1.54 ;
      RECT  13.38 1.54 13.715 1.545 ;
      RECT  13.385 1.545 13.72 1.55 ;
      RECT  13.39 1.55 13.725 1.555 ;
      RECT  13.395 1.555 13.73 1.56 ;
      RECT  13.4 1.56 13.735 1.565 ;
      RECT  13.405 1.565 16.915 1.57 ;
      RECT  13.41 1.57 16.915 1.575 ;
      RECT  13.415 1.575 16.915 1.58 ;
      RECT  13.42 1.58 16.915 1.585 ;
      RECT  13.425 1.585 16.915 1.59 ;
      RECT  13.43 1.59 16.915 1.595 ;
      RECT  13.435 1.595 16.915 1.6 ;
      RECT  13.44 1.6 16.915 1.605 ;
      RECT  13.445 1.605 16.915 1.61 ;
      RECT  13.45 1.61 16.915 1.615 ;
      RECT  13.455 1.615 16.915 1.62 ;
      RECT  13.46 1.62 16.915 1.625 ;
      RECT  13.465 1.625 16.915 1.63 ;
      RECT  13.47 1.63 16.915 1.635 ;
      RECT  13.475 1.635 16.915 1.64 ;
      RECT  13.48 1.64 16.915 1.645 ;
      RECT  13.485 1.645 16.915 1.65 ;
      RECT  13.49 1.65 16.915 1.655 ;
      RECT  13.495 1.655 16.915 1.66 ;
      RECT  13.5 1.66 16.915 1.665 ;
      RECT  13.505 1.665 16.915 1.67 ;
      RECT  13.51 1.67 16.915 1.675 ;
      RECT  13.515 1.675 16.915 1.68 ;
      RECT  13.52 1.68 16.915 1.685 ;
      RECT  13.525 1.685 16.915 1.69 ;
      RECT  13.53 1.69 16.915 1.695 ;
      RECT  13.535 1.695 16.915 1.7 ;
      RECT  13.54 1.7 16.915 1.705 ;
      RECT  13.545 1.705 16.915 1.71 ;
      RECT  13.55 1.71 16.915 1.715 ;
      RECT  13.555 1.715 16.915 1.72 ;
      RECT  13.56 1.72 16.915 1.725 ;
      RECT  13.565 1.725 16.915 1.73 ;
      RECT  13.57 1.73 16.915 1.735 ;
      RECT  13.575 1.735 16.915 1.74 ;
      RECT  13.58 1.74 16.915 1.745 ;
      RECT  13.585 1.745 16.915 1.75 ;
      RECT  13.59 1.75 16.915 1.755 ;
      RECT  13.595 1.755 16.915 1.76 ;
      RECT  13.6 1.76 16.915 1.765 ;
      RECT  13.605 1.765 16.915 1.77 ;
      RECT  13.61 1.77 16.915 1.775 ;
      RECT  13.615 1.775 16.915 1.78 ;
      RECT  13.62 1.78 16.915 1.785 ;
      RECT  13.625 1.785 16.915 1.79 ;
      RECT  13.63 1.79 16.915 1.795 ;
      RECT  17.4 1.565 18.595 1.795 ;
      RECT  18.365 1.795 18.595 2.405 ;
      RECT  18.365 2.405 22.01 2.635 ;
      RECT  18.365 2.635 18.595 3.245 ;
      RECT  15.86 3.245 18.595 3.475 ;
      RECT  23.965 1.565 24.46 1.795 ;
      RECT  23.965 1.795 24.195 2.405 ;
      RECT  23.965 2.405 26.49 2.635 ;
      RECT  23.965 2.635 24.195 3.245 ;
      RECT  23.965 3.245 24.46 3.475 ;
      RECT  6.2 1.75 6.835 1.98 ;
      RECT  6.605 1.98 6.835 2.405 ;
      RECT  6.605 2.405 7.45 2.635 ;
      RECT  6.605 2.635 6.835 3.16 ;
      RECT  6.2 3.16 6.835 3.39 ;
      RECT  7.67 1.75 8.01 1.98 ;
      RECT  7.725 1.98 7.955 2.685 ;
      RECT  7.725 2.685 9.175 2.915 ;
      RECT  8.795 2.66 9.175 2.685 ;
      RECT  8.795 2.915 9.175 2.94 ;
      RECT  7.725 2.915 7.955 3.315 ;
      RECT  9.14 1.75 10.095 1.98 ;
      RECT  9.865 1.98 10.095 3.68 ;
      RECT  8.585 3.68 10.095 3.91 ;
      RECT  8.585 3.91 8.815 4.02 ;
      RECT  7.725 4.02 8.815 4.25 ;
      RECT  7.725 4.25 7.955 4.54 ;
      RECT  4.925 4.54 7.955 4.77 ;
      RECT  4.925 4.77 5.155 5.0 ;
      RECT  3.75 5.0 5.155 5.23 ;
      RECT  12.15 1.75 12.49 1.98 ;
      RECT  12.205 1.98 12.435 3.315 ;
      RECT  12.765 1.75 13.26 1.98 ;
      RECT  12.765 1.98 12.995 2.445 ;
      RECT  12.765 2.445 14.17 2.675 ;
      RECT  12.765 2.675 12.995 3.32 ;
      RECT  12.76 3.32 12.995 3.325 ;
      RECT  12.755 3.325 12.995 3.33 ;
      RECT  12.75 3.33 12.995 3.335 ;
      RECT  12.745 3.335 12.995 3.34 ;
      RECT  12.74 3.34 12.995 3.345 ;
      RECT  12.735 3.345 12.995 3.35 ;
      RECT  12.73 3.35 12.995 3.355 ;
      RECT  12.725 3.355 12.995 3.36 ;
      RECT  12.72 3.36 12.995 3.365 ;
      RECT  12.715 3.365 12.995 3.37 ;
      RECT  12.71 3.37 12.995 3.375 ;
      RECT  12.705 3.375 12.995 3.38 ;
      RECT  12.7 3.38 12.995 3.385 ;
      RECT  12.695 3.385 12.995 3.39 ;
      RECT  12.69 3.39 12.995 3.395 ;
      RECT  12.685 3.395 12.995 3.4 ;
      RECT  12.68 3.4 12.995 3.405 ;
      RECT  12.675 3.405 12.995 3.41 ;
      RECT  12.67 3.41 12.995 3.415 ;
      RECT  12.665 3.415 12.99 3.42 ;
      RECT  12.66 3.42 12.985 3.425 ;
      RECT  12.655 3.425 12.98 3.43 ;
      RECT  12.65 3.43 12.975 3.435 ;
      RECT  12.645 3.435 12.97 3.44 ;
      RECT  12.64 3.44 12.965 3.445 ;
      RECT  12.635 3.445 12.96 3.45 ;
      RECT  12.63 3.45 12.955 3.455 ;
      RECT  12.625 3.455 12.95 3.46 ;
      RECT  12.62 3.46 12.945 3.465 ;
      RECT  12.615 3.465 12.94 3.47 ;
      RECT  12.61 3.47 12.935 3.475 ;
      RECT  12.605 3.475 12.93 3.48 ;
      RECT  12.6 3.48 12.925 3.485 ;
      RECT  12.595 3.485 12.92 3.49 ;
      RECT  12.59 3.49 12.915 3.495 ;
      RECT  12.585 3.495 12.91 3.5 ;
      RECT  12.58 3.5 12.905 3.505 ;
      RECT  12.575 3.505 12.9 3.51 ;
      RECT  12.57 3.51 12.895 3.515 ;
      RECT  12.565 3.515 12.89 3.52 ;
      RECT  12.56 3.52 12.885 3.525 ;
      RECT  12.555 3.525 12.88 3.53 ;
      RECT  12.55 3.53 12.875 3.535 ;
      RECT  12.545 3.535 12.87 3.54 ;
      RECT  12.54 3.54 12.865 3.545 ;
      RECT  12.535 3.545 12.86 3.55 ;
      RECT  12.53 3.55 12.855 3.555 ;
      RECT  10.68 1.75 11.315 1.98 ;
      RECT  11.085 1.98 11.315 3.555 ;
      RECT  10.68 3.555 12.85 3.56 ;
      RECT  10.68 3.56 12.845 3.565 ;
      RECT  10.68 3.565 12.84 3.57 ;
      RECT  10.68 3.57 12.835 3.575 ;
      RECT  10.68 3.575 12.83 3.58 ;
      RECT  10.68 3.58 12.825 3.585 ;
      RECT  10.68 3.585 12.82 3.59 ;
      RECT  10.68 3.59 12.815 3.595 ;
      RECT  10.68 3.595 12.81 3.6 ;
      RECT  10.68 3.6 12.805 3.605 ;
      RECT  10.68 3.605 12.8 3.61 ;
      RECT  10.68 3.61 12.795 3.615 ;
      RECT  10.68 3.615 12.79 3.62 ;
      RECT  10.68 3.62 12.785 3.625 ;
      RECT  10.68 3.625 12.78 3.63 ;
      RECT  10.68 3.63 12.775 3.635 ;
      RECT  10.68 3.635 12.77 3.64 ;
      RECT  10.68 3.64 12.765 3.645 ;
      RECT  10.68 3.645 12.76 3.65 ;
      RECT  10.68 3.65 12.755 3.655 ;
      RECT  10.68 3.655 12.75 3.66 ;
      RECT  10.68 3.66 12.745 3.665 ;
      RECT  10.68 3.665 12.74 3.67 ;
      RECT  10.68 3.67 12.735 3.675 ;
      RECT  10.68 3.675 12.73 3.68 ;
      RECT  10.68 3.68 12.725 3.685 ;
      RECT  10.68 3.685 12.72 3.69 ;
      RECT  10.68 3.69 12.715 3.695 ;
      RECT  10.68 3.695 12.71 3.7 ;
      RECT  10.68 3.7 12.705 3.705 ;
      RECT  10.68 3.705 12.7 3.71 ;
      RECT  10.68 3.71 12.695 3.715 ;
      RECT  10.68 3.715 12.69 3.72 ;
      RECT  10.68 3.72 12.685 3.725 ;
      RECT  10.68 3.725 12.68 3.73 ;
      RECT  10.68 3.73 12.675 3.735 ;
      RECT  10.68 3.735 12.67 3.74 ;
      RECT  10.68 3.74 12.665 3.745 ;
      RECT  10.68 3.745 12.66 3.75 ;
      RECT  10.68 3.75 12.655 3.755 ;
      RECT  10.68 3.755 12.65 3.76 ;
      RECT  10.68 3.76 12.645 3.765 ;
      RECT  10.68 3.765 12.64 3.77 ;
      RECT  10.68 3.77 12.635 3.775 ;
      RECT  10.68 3.775 12.63 3.78 ;
      RECT  10.68 3.78 12.625 3.785 ;
      RECT  27.27 2.405 28.73 2.635 ;
      RECT  5.485 2.41 6.33 2.64 ;
      RECT  5.485 2.64 5.715 3.16 ;
      RECT  4.66 3.16 5.715 3.39 ;
      RECT  10.525 2.21 10.755 2.66 ;
      RECT  10.325 2.66 10.755 2.94 ;
      RECT  9.405 2.35 9.635 3.22 ;
      RECT  8.385 3.22 9.635 3.225 ;
      RECT  8.38 3.225 9.635 3.23 ;
      RECT  8.375 3.23 9.635 3.235 ;
      RECT  8.37 3.235 9.635 3.24 ;
      RECT  8.365 3.24 9.635 3.245 ;
      RECT  8.36 3.245 9.635 3.25 ;
      RECT  8.355 3.25 9.635 3.255 ;
      RECT  8.35 3.255 9.635 3.26 ;
      RECT  8.345 3.26 9.635 3.265 ;
      RECT  8.34 3.265 9.635 3.27 ;
      RECT  8.335 3.27 9.635 3.275 ;
      RECT  8.33 3.275 9.635 3.28 ;
      RECT  8.325 3.28 9.635 3.285 ;
      RECT  8.32 3.285 9.635 3.29 ;
      RECT  8.315 3.29 9.635 3.295 ;
      RECT  8.31 3.295 9.635 3.3 ;
      RECT  8.305 3.3 9.635 3.305 ;
      RECT  8.3 3.305 9.635 3.31 ;
      RECT  8.295 3.31 9.635 3.315 ;
      RECT  8.29 3.315 9.635 3.32 ;
      RECT  8.285 3.32 9.635 3.325 ;
      RECT  8.28 3.325 9.635 3.33 ;
      RECT  8.275 3.33 9.635 3.335 ;
      RECT  8.27 3.335 9.635 3.34 ;
      RECT  8.265 3.34 9.635 3.345 ;
      RECT  8.26 3.345 9.635 3.35 ;
      RECT  8.255 3.35 9.635 3.355 ;
      RECT  8.25 3.355 9.635 3.36 ;
      RECT  8.245 3.36 9.635 3.365 ;
      RECT  8.24 3.365 9.635 3.37 ;
      RECT  8.235 3.37 9.635 3.375 ;
      RECT  8.23 3.375 9.635 3.38 ;
      RECT  8.225 3.38 9.635 3.385 ;
      RECT  8.22 3.385 9.635 3.39 ;
      RECT  8.215 3.39 9.635 3.395 ;
      RECT  8.21 3.395 9.635 3.4 ;
      RECT  8.205 3.4 9.635 3.405 ;
      RECT  8.2 3.405 9.635 3.41 ;
      RECT  8.195 3.41 9.635 3.415 ;
      RECT  8.19 3.415 9.635 3.42 ;
      RECT  8.185 3.42 9.635 3.425 ;
      RECT  8.18 3.425 9.635 3.43 ;
      RECT  8.175 3.43 9.635 3.435 ;
      RECT  8.17 3.435 9.635 3.44 ;
      RECT  8.165 3.44 9.635 3.445 ;
      RECT  8.16 3.445 9.635 3.45 ;
      RECT  8.155 3.45 8.48 3.455 ;
      RECT  8.15 3.455 8.475 3.46 ;
      RECT  8.145 3.46 8.47 3.465 ;
      RECT  8.14 3.465 8.465 3.47 ;
      RECT  8.135 3.47 8.46 3.475 ;
      RECT  8.13 3.475 8.455 3.48 ;
      RECT  8.125 3.48 8.45 3.485 ;
      RECT  8.12 3.485 8.445 3.49 ;
      RECT  8.115 3.49 8.44 3.495 ;
      RECT  8.11 3.495 8.435 3.5 ;
      RECT  8.105 3.5 8.43 3.505 ;
      RECT  8.1 3.505 8.425 3.51 ;
      RECT  8.095 3.51 8.42 3.515 ;
      RECT  8.09 3.515 8.415 3.52 ;
      RECT  8.085 3.52 8.41 3.525 ;
      RECT  8.08 3.525 8.405 3.53 ;
      RECT  8.075 3.53 8.4 3.535 ;
      RECT  8.07 3.535 8.395 3.54 ;
      RECT  8.065 3.54 8.39 3.545 ;
      RECT  8.06 3.545 8.385 3.55 ;
      RECT  8.055 3.55 8.38 3.555 ;
      RECT  8.05 3.555 8.375 3.56 ;
      RECT  7.165 3.56 8.37 3.565 ;
      RECT  7.165 3.565 8.365 3.57 ;
      RECT  7.165 3.57 8.36 3.575 ;
      RECT  7.165 3.575 8.355 3.58 ;
      RECT  7.165 3.58 8.35 3.585 ;
      RECT  7.165 3.585 8.345 3.59 ;
      RECT  7.165 3.59 8.34 3.595 ;
      RECT  7.165 3.595 8.335 3.6 ;
      RECT  7.165 3.6 8.33 3.605 ;
      RECT  7.165 3.605 8.325 3.61 ;
      RECT  7.165 3.61 8.32 3.615 ;
      RECT  7.165 3.615 8.315 3.62 ;
      RECT  3.805 3.62 8.31 3.625 ;
      RECT  3.805 3.625 8.305 3.63 ;
      RECT  3.805 3.63 8.3 3.635 ;
      RECT  3.805 3.635 8.295 3.64 ;
      RECT  3.805 3.64 8.29 3.645 ;
      RECT  3.805 3.645 8.285 3.65 ;
      RECT  3.805 3.65 8.28 3.655 ;
      RECT  3.805 3.655 8.275 3.66 ;
      RECT  3.805 3.66 8.27 3.665 ;
      RECT  3.805 3.665 8.265 3.67 ;
      RECT  3.805 3.67 8.26 3.675 ;
      RECT  3.805 3.675 8.255 3.68 ;
      RECT  3.805 3.68 8.25 3.685 ;
      RECT  3.805 3.685 8.245 3.69 ;
      RECT  3.805 3.69 8.24 3.695 ;
      RECT  3.805 3.695 8.235 3.7 ;
      RECT  3.805 3.7 8.23 3.705 ;
      RECT  3.805 3.705 8.225 3.71 ;
      RECT  3.805 3.71 8.22 3.715 ;
      RECT  3.805 3.715 8.215 3.72 ;
      RECT  3.805 3.72 8.21 3.725 ;
      RECT  3.805 3.725 8.205 3.73 ;
      RECT  3.805 3.73 8.2 3.735 ;
      RECT  3.805 3.735 8.195 3.74 ;
      RECT  3.805 3.74 8.19 3.745 ;
      RECT  3.805 3.745 8.185 3.75 ;
      RECT  3.805 3.75 8.18 3.755 ;
      RECT  3.805 3.755 8.175 3.76 ;
      RECT  3.805 3.76 8.17 3.765 ;
      RECT  3.805 3.765 8.165 3.77 ;
      RECT  3.805 3.77 8.16 3.775 ;
      RECT  3.805 3.775 8.155 3.78 ;
      RECT  3.805 3.78 8.15 3.785 ;
      RECT  3.805 3.785 8.145 3.79 ;
      RECT  3.805 3.79 7.395 3.85 ;
      RECT  3.805 3.85 4.035 4.08 ;
      RECT  2.685 4.08 4.035 4.31 ;
      RECT  2.685 4.31 2.915 5.0 ;
      RECT  1.51 5.0 2.915 5.23 ;
      RECT  1.72 3.16 2.76 3.39 ;
      RECT  3.245 3.16 4.3 3.39 ;
      RECT  3.245 3.39 3.475 3.62 ;
      RECT  2.125 3.62 3.475 3.85 ;
      RECT  2.125 3.85 2.355 4.365 ;
      RECT  0.18 4.365 2.355 4.595 ;
      RECT  13.065 3.7 15.5 3.93 ;
      RECT  13.065 3.93 13.295 4.015 ;
      RECT  12.205 4.015 13.295 4.145 ;
      RECT  9.045 4.145 13.295 4.245 ;
      RECT  9.045 4.245 12.435 4.375 ;
      RECT  9.045 4.375 9.275 4.48 ;
      RECT  8.44 4.48 9.275 4.71 ;
      RECT  15.73 3.805 18.44 4.035 ;
      RECT  15.73 4.035 15.96 4.16 ;
      RECT  13.525 4.16 15.96 4.39 ;
      RECT  13.525 4.39 13.755 4.475 ;
      RECT  12.92 4.475 13.755 4.705 ;
      RECT  4.365 4.08 7.24 4.31 ;
      RECT  4.365 4.31 4.595 4.54 ;
      RECT  3.19 4.54 4.595 4.77 ;
      RECT  16.19 4.365 17.42 4.595 ;
      RECT  16.19 4.595 16.42 4.62 ;
      RECT  17.19 4.595 17.42 5.0 ;
      RECT  13.985 4.62 16.42 4.85 ;
      RECT  13.985 4.85 14.215 4.935 ;
      RECT  12.15 4.935 14.215 5.165 ;
      RECT  17.19 5.0 17.53 5.23 ;
      RECT  9.505 4.61 10.755 4.84 ;
      RECT  9.505 4.84 9.735 5.0 ;
      RECT  10.525 4.84 10.755 5.0 ;
      RECT  5.99 5.0 9.735 5.23 ;
      RECT  10.525 5.0 11.92 5.23 ;
      LAYER METAL2 ;
      RECT  8.795 2.66 10.755 2.94 ;
      LAYER VIA12 ;
      RECT  8.855 2.67 9.115 2.93 ;
      RECT  10.435 2.67 10.695 2.93 ;
  END
END MDN_FSDPRB_4